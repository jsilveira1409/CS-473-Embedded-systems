// DE0_Nano_SOPC.v

// Generated using ACDS version 13.1 162 at 2014.07.02.13:44:20

`timescale 1 ps / 1 ps
module DE0_Nano_SOPC (
		input  wire [1:0]  in_port_to_the_key,                               //                   key_external_connection.export
		input  wire        clk_50,                                           //                             clk_50_clk_in.clk
		output wire        locked_from_the_altpll_sys,                       //                 altpll_sys_locked_conduit.export
		input  wire        reset_n,                                          //                       clk_50_clk_in_reset.reset_n
		output wire [7:0]  out_port_from_the_led,                            //                   led_external_connection.export
		output wire        phasedone_from_the_altpll_sys,                    //              altpll_sys_phasedone_conduit.export
		output wire [12:0] zs_addr_from_the_sdram,                           //                                sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                             //                                          .ba
		output wire        zs_cas_n_from_the_sdram,                          //                                          .cas_n
		output wire        zs_cke_from_the_sdram,                            //                                          .cke
		output wire        zs_cs_n_from_the_sdram,                           //                                          .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram,                      //                                          .dq
		output wire [1:0]  zs_dqm_from_the_sdram,                            //                                          .dqm
		output wire        zs_ras_n_from_the_sdram,                          //                                          .ras_n
		output wire        zs_we_n_from_the_sdram,                           //                                          .we_n
		input  wire [3:0]  in_port_to_the_sw,                                //                    sw_external_connection.export
		output wire        altpll_sys_c3_out,                                //                             altpll_sys_c3.clk
		output wire        altpll_sdram,                                     //                             altpll_sys_c1.clk
		output wire        lt24_controller_0_conduit_end_cs,                 //             lt24_controller_0_conduit_end.cs
		output wire        lt24_controller_0_conduit_end_rs,                 //                                          .rs
		output wire        lt24_controller_0_conduit_end_rd,                 //                                          .rd
		output wire        lt24_controller_0_conduit_end_wr,                 //                                          .wr
		output wire [15:0] lt24_controller_0_conduit_end_data,               //                                          .data
		output wire        lcd_reset_n_external_connection_export,           //           lcd_reset_n_external_connection.export
		input  wire        touch_panel_spi_external_MISO,                    //                  touch_panel_spi_external.MISO
		output wire        touch_panel_spi_external_MOSI,                    //                                          .MOSI
		output wire        touch_panel_spi_external_SCLK,                    //                                          .SCLK
		output wire        touch_panel_spi_external_SS_n,                    //                                          .SS_n
		input  wire        touch_panel_pen_irq_n_external_connection_export, // touch_panel_pen_irq_n_external_connection.export
		input  wire        touch_panel_busy_external_connection_export,      //      touch_panel_busy_external_connection.export
		output wire        epcs_flash_controller_0_external_dclk,            //          epcs_flash_controller_0_external.dclk
		output wire        epcs_flash_controller_0_external_sce,             //                                          .sce
		output wire        epcs_flash_controller_0_external_sdo,             //                                          .sdo
		input  wire        epcs_flash_controller_0_external_data0            //                                          .data0
	);

	wire         altpll_sys_c0_clk;                                                      // altpll_sys:c0 -> [LCD_RESET_N:clk, LT24_Controller_0:clk, clock_crossing_io:s0_clk, cpu:clk, epcs_flash_controller_0:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, jtag_uart:clk, mm_interconnect_0:altpll_sys_c0_clk, rst_controller_002:clk, sdram:clk, touch_panel_busy:clk, touch_panel_pen_irq_n:clk, touch_panel_spi:clk]
	wire         altpll_sys_c2_clk;                                                      // altpll_sys:c2 -> [clock_crossing_io:m0_clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, key:clk, led:clk, mm_interconnect_1:altpll_sys_c2_clk, rst_controller:clk, sw:clk, sysid:clock, timer:clk]
	wire         cpu_jtag_debug_module_reset_reset;                                      // cpu:jtag_debug_module_resetrequest -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, sdram:reset_n]
	wire  [31:0] mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata;           // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_writedata -> LT24_Controller_0:s_writedata
	wire   [0:0] mm_interconnect_0_lt24_controller_0_avalon_slave_0_address;             // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_address -> LT24_Controller_0:s_address
	wire         mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect;          // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_chipselect -> LT24_Controller_0:s_chipselect_n
	wire         mm_interconnect_0_lt24_controller_0_avalon_slave_0_write;               // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_write -> LT24_Controller_0:s_write_n
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_writedata;           // mm_interconnect_0:touch_panel_spi_spi_control_port_writedata -> touch_panel_spi:data_from_cpu
	wire   [2:0] mm_interconnect_0_touch_panel_spi_spi_control_port_address;             // mm_interconnect_0:touch_panel_spi_spi_control_port_address -> touch_panel_spi:mem_addr
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect;          // mm_interconnect_0:touch_panel_spi_spi_control_port_chipselect -> touch_panel_spi:spi_select
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_write;               // mm_interconnect_0:touch_panel_spi_spi_control_port_write -> touch_panel_spi:write_n
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_read;                // mm_interconnect_0:touch_panel_spi_spi_control_port_read -> touch_panel_spi:read_n
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_readdata;            // touch_panel_spi:data_to_cpu -> mm_interconnect_0:touch_panel_spi_spi_control_port_readdata
	wire   [1:0] mm_interconnect_0_touch_panel_busy_s1_address;                          // mm_interconnect_0:touch_panel_busy_s1_address -> touch_panel_busy:address
	wire  [31:0] mm_interconnect_0_touch_panel_busy_s1_readdata;                         // touch_panel_busy:readdata -> mm_interconnect_0:touch_panel_busy_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;              // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                 // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         cpu_instruction_master_waitrequest;                                     // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                         // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                            // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                        // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                                   // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;                       // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire   [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;                         // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire         mm_interconnect_0_altpll_sys_pll_slave_write;                           // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire         mm_interconnect_0_altpll_sys_pll_slave_read;                            // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;                        // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire  [31:0] mm_interconnect_0_lcd_reset_n_s1_writedata;                             // mm_interconnect_0:LCD_RESET_N_s1_writedata -> LCD_RESET_N:writedata
	wire   [1:0] mm_interconnect_0_lcd_reset_n_s1_address;                               // mm_interconnect_0:LCD_RESET_N_s1_address -> LCD_RESET_N:address
	wire         mm_interconnect_0_lcd_reset_n_s1_chipselect;                            // mm_interconnect_0:LCD_RESET_N_s1_chipselect -> LCD_RESET_N:chipselect
	wire         mm_interconnect_0_lcd_reset_n_s1_write;                                 // mm_interconnect_0:LCD_RESET_N_s1_write -> LCD_RESET_N:write_n
	wire  [31:0] mm_interconnect_0_lcd_reset_n_s1_readdata;                              // LCD_RESET_N:readdata -> mm_interconnect_0:LCD_RESET_N_s1_readdata
	wire  [31:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata;                   // mm_interconnect_0:touch_panel_pen_irq_n_s1_writedata -> touch_panel_pen_irq_n:writedata
	wire   [1:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_address;                     // mm_interconnect_0:touch_panel_pen_irq_n_s1_address -> touch_panel_pen_irq_n:address
	wire         mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect;                  // mm_interconnect_0:touch_panel_pen_irq_n_s1_chipselect -> touch_panel_pen_irq_n:chipselect
	wire         mm_interconnect_0_touch_panel_pen_irq_n_s1_write;                       // mm_interconnect_0:touch_panel_pen_irq_n_s1_write -> touch_panel_pen_irq_n:write_n
	wire  [31:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata;                    // touch_panel_pen_irq_n:readdata -> mm_interconnect_0:touch_panel_pen_irq_n_s1_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                     // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                      // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                       // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [6:0] mm_interconnect_0_clock_crossing_io_s0_address;                         // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                           // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                            // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                        // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                     // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                   // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                      // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                    // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                      // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                        // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                          // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                           // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                       // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                    // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                     // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_writedata -> epcs_flash_controller_0:writedata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_address -> epcs_flash_controller_0:address
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_chipselect -> epcs_flash_controller_0:chipselect
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_write -> epcs_flash_controller_0:write_n
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_read -> epcs_flash_controller_0:read_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata;   // epcs_flash_controller_0:readdata -> mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_readdata
	wire         cpu_data_master_waitrequest;                                            // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                              // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [26:0] cpu_data_master_address;                                                // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                                  // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                                   // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                               // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                            // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire         cpu_data_master_readdatavalid;                                          // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                             // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                 // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                   // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                     // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                  // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                       // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                        // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                    // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                               // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                  // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                                      // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                        // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_chipselect;                                     // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire         mm_interconnect_1_sw_s1_write;                                          // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                       // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                          // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                         // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                     // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                       // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_chipselect;                                    // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire         mm_interconnect_1_key_s1_write;                                         // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                      // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [0:0] clock_crossing_io_m0_burstcount;                                        // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire         clock_crossing_io_m0_waitrequest;                                       // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire   [6:0] clock_crossing_io_m0_address;                                           // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire  [31:0] clock_crossing_io_m0_writedata;                                         // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                             // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire         clock_crossing_io_m0_read;                                              // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire  [31:0] clock_crossing_io_m0_readdata;                                          // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                       // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [3:0] clock_crossing_io_m0_byteenable;                                        // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                     // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                                   // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                                     // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_chipselect;                                  // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_1_timer_s1_write;                                       // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                                    // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                     // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                       // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_chipselect;                                    // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_1_led_s1_write;                                         // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                      // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire         irq_mapper_receiver3_irq;                                               // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                               // touch_panel_spi:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                               // touch_panel_pen_irq_n:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                               // epcs_flash_controller_0:irq -> irq_mapper:receiver6_irq
	wire  [31:0] cpu_d_irq_irq;                                                          // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                               // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                          // timer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                               // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                      // key:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                               // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                      // sw:irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [clock_crossing_io:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, key:reset_n, led:reset_n, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, sw:reset_n, sysid:reset_n, timer:reset_n]
	wire         rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> [altpll_sys:reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                     // rst_controller_002:reset_out -> [LCD_RESET_N:reset_n, LT24_Controller_0:reset_n, clock_crossing_io:s0_reset, cpu:reset_n, epcs_flash_controller_0:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, touch_panel_busy:reset_n, touch_panel_pen_irq_n:reset_n, touch_panel_spi:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                                 // rst_controller_002:reset_req -> [cpu:reset_req, epcs_flash_controller_0:reset_req, rst_translator:reset_req_in]

	DE0_Nano_SOPC_timer timer (
		.clk        (altpll_sys_c2_clk),                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	DE0_Nano_SOPC_key key (
		.clk        (altpll_sys_c2_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_key),                  // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)    //                 irq.irq
	);

	DE0_Nano_SOPC_sw sw (
		.clk        (altpll_sys_c2_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_sw),                  // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)   //                 irq.irq
	);

	DE0_Nano_SOPC_led led (
		.clk        (altpll_sys_c2_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led)                // external_connection.export
	);

	DE0_Nano_SOPC_sdram sdram (
		.clk            (altpll_sys_c0_clk),                        //   clk.clk
		.reset_n        (~cpu_jtag_debug_module_reset_reset),       // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	DE0_Nano_SOPC_altpll_sys altpll_sys (
		.clk       (clk_50),                                           //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0        (altpll_sys_c0_clk),                                //                    c0.clk
		.c1        (altpll_sdram),                                     //                    c1.clk
		.c2        (altpll_sys_c2_clk),                                //                    c2.clk
		.c3        (altpll_sys_c3_out),                                //                    c3.clk
		.c4        (),                                                 //                    c4.clk
		.areset    (),                                                 //        areset_conduit.export
		.locked    (locked_from_the_altpll_sys),                       //        locked_conduit.export
		.phasedone (phasedone_from_the_altpll_sys)                     //     phasedone_conduit.export
	);

	DE0_Nano_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_sys_c0_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (7),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_sys_c2_clk),                                    //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (altpll_sys_c0_clk),                                    //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE0_Nano_SOPC_cpu cpu (
		.clk                                   (altpll_sys_c0_clk),                                   //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE0_Nano_SOPC_sysid sysid (
		.clock    (altpll_sys_c2_clk),                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	LT24_Controller lt24_controller_0 (
		.clk            (altpll_sys_c0_clk),                                              //          clock.clk
		.reset_n        (~rst_controller_002_reset_out_reset),                            //          reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect_n
		.s_write_n      (~mm_interconnect_0_lt24_controller_0_avalon_slave_0_write),      //               .write_n
		.s_writedata    (mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata),   //               .writedata
		.s_address      (mm_interconnect_0_lt24_controller_0_avalon_slave_0_address),     //               .address
		.lt24_cs        (lt24_controller_0_conduit_end_cs),                               //    conduit_end.export
		.lt24_rs        (lt24_controller_0_conduit_end_rs),                               //               .export
		.lt24_rd        (lt24_controller_0_conduit_end_rd),                               //               .export
		.lt24_wr        (lt24_controller_0_conduit_end_wr),                               //               .export
		.lt24_data      (lt24_controller_0_conduit_end_data)                              //               .export
	);

	DE0_Nano_SOPC_LCD_RESET_N lcd_reset_n (
		.clk        (altpll_sys_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_lcd_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_reset_n_s1_readdata),   //                    .readdata
		.out_port   (lcd_reset_n_external_connection_export)       // external_connection.export
	);

	DE0_Nano_SOPC_touch_panel_pen_irq_n touch_panel_pen_irq_n (
		.clk        (altpll_sys_c0_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_touch_panel_pen_irq_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_panel_pen_irq_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata),   //                    .readdata
		.in_port    (touch_panel_pen_irq_n_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                               //                 irq.irq
	);

	DE0_Nano_SOPC_touch_panel_busy touch_panel_busy (
		.clk      (altpll_sys_c0_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_touch_panel_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touch_panel_busy_s1_readdata), //                    .readdata
		.in_port  (touch_panel_busy_external_connection_export)     // external_connection.export
	);

	DE0_Nano_SOPC_touch_panel_spi touch_panel_spi (
		.clk           (altpll_sys_c0_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                           //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_touch_panel_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_touch_panel_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver4_irq),                                      //              irq.irq
		.MISO          (touch_panel_spi_external_MISO),                                 //         external.export
		.MOSI          (touch_panel_spi_external_MOSI),                                 //                 .export
		.SCLK          (touch_panel_spi_external_SCLK),                                 //                 .export
		.SS_n          (touch_panel_spi_external_SS_n)                                  //                 .export
	);

	DE0_Nano_SOPC_epcs_flash_controller_0 epcs_flash_controller_0 (
		.clk           (altpll_sys_c0_clk),                                                      //               clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                                    //             reset.reset_n
		.reset_req     (rst_controller_002_reset_out_reset_req),                                 //                  .reset_req
		.address       (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                                       //                  .dataavailable
		.endofpacket   (),                                                                       //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                                       //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver6_irq),                                               //               irq.irq
		.dclk          (epcs_flash_controller_0_external_dclk),                                  //          external.export
		.sce           (epcs_flash_controller_0_external_sce),                                   //                  .export
		.sdo           (epcs_flash_controller_0_external_sdo),                                   //                  .export
		.data0         (epcs_flash_controller_0_external_data0)                                  //                  .export
	);

	DE0_Nano_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c0_clk                                            (altpll_sys_c0_clk),                                                      //                                          altpll_sys_c0.clk
		.clk_50_clk_clk                                               (clk_50),                                                                 //                                             clk_50_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                     // altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                      (rst_controller_002_reset_out_reset),                                     //                      cpu_reset_n_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset                      (cpu_jtag_debug_module_reset_reset),                                      //                      sdram_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                      (cpu_data_master_address),                                                //                                        cpu_data_master.address
		.cpu_data_master_waitrequest                                  (cpu_data_master_waitrequest),                                            //                                                       .waitrequest
		.cpu_data_master_byteenable                                   (cpu_data_master_byteenable),                                             //                                                       .byteenable
		.cpu_data_master_read                                         (cpu_data_master_read),                                                   //                                                       .read
		.cpu_data_master_readdata                                     (cpu_data_master_readdata),                                               //                                                       .readdata
		.cpu_data_master_readdatavalid                                (cpu_data_master_readdatavalid),                                          //                                                       .readdatavalid
		.cpu_data_master_write                                        (cpu_data_master_write),                                                  //                                                       .write
		.cpu_data_master_writedata                                    (cpu_data_master_writedata),                                              //                                                       .writedata
		.cpu_data_master_debugaccess                                  (cpu_data_master_debugaccess),                                            //                                                       .debugaccess
		.cpu_instruction_master_address                               (cpu_instruction_master_address),                                         //                                 cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                           (cpu_instruction_master_waitrequest),                                     //                                                       .waitrequest
		.cpu_instruction_master_read                                  (cpu_instruction_master_read),                                            //                                                       .read
		.cpu_instruction_master_readdata                              (cpu_instruction_master_readdata),                                        //                                                       .readdata
		.cpu_instruction_master_readdatavalid                         (cpu_instruction_master_readdatavalid),                                   //                                                       .readdatavalid
		.altpll_sys_pll_slave_address                                 (mm_interconnect_0_altpll_sys_pll_slave_address),                         //                                   altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                   (mm_interconnect_0_altpll_sys_pll_slave_write),                           //                                                       .write
		.altpll_sys_pll_slave_read                                    (mm_interconnect_0_altpll_sys_pll_slave_read),                            //                                                       .read
		.altpll_sys_pll_slave_readdata                                (mm_interconnect_0_altpll_sys_pll_slave_readdata),                        //                                                       .readdata
		.altpll_sys_pll_slave_writedata                               (mm_interconnect_0_altpll_sys_pll_slave_writedata),                       //                                                       .writedata
		.clock_crossing_io_s0_address                                 (mm_interconnect_0_clock_crossing_io_s0_address),                         //                                   clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                                   (mm_interconnect_0_clock_crossing_io_s0_write),                           //                                                       .write
		.clock_crossing_io_s0_read                                    (mm_interconnect_0_clock_crossing_io_s0_read),                            //                                                       .read
		.clock_crossing_io_s0_readdata                                (mm_interconnect_0_clock_crossing_io_s0_readdata),                        //                                                       .readdata
		.clock_crossing_io_s0_writedata                               (mm_interconnect_0_clock_crossing_io_s0_writedata),                       //                                                       .writedata
		.clock_crossing_io_s0_burstcount                              (mm_interconnect_0_clock_crossing_io_s0_burstcount),                      //                                                       .burstcount
		.clock_crossing_io_s0_byteenable                              (mm_interconnect_0_clock_crossing_io_s0_byteenable),                      //                                                       .byteenable
		.clock_crossing_io_s0_readdatavalid                           (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),                   //                                                       .readdatavalid
		.clock_crossing_io_s0_waitrequest                             (mm_interconnect_0_clock_crossing_io_s0_waitrequest),                     //                                                       .waitrequest
		.clock_crossing_io_s0_debugaccess                             (mm_interconnect_0_clock_crossing_io_s0_debugaccess),                     //                                                       .debugaccess
		.cpu_jtag_debug_module_address                                (mm_interconnect_0_cpu_jtag_debug_module_address),                        //                                  cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                                  (mm_interconnect_0_cpu_jtag_debug_module_write),                          //                                                       .write
		.cpu_jtag_debug_module_read                                   (mm_interconnect_0_cpu_jtag_debug_module_read),                           //                                                       .read
		.cpu_jtag_debug_module_readdata                               (mm_interconnect_0_cpu_jtag_debug_module_readdata),                       //                                                       .readdata
		.cpu_jtag_debug_module_writedata                              (mm_interconnect_0_cpu_jtag_debug_module_writedata),                      //                                                       .writedata
		.cpu_jtag_debug_module_byteenable                             (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                     //                                                       .byteenable
		.cpu_jtag_debug_module_waitrequest                            (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                    //                                                       .waitrequest
		.cpu_jtag_debug_module_debugaccess                            (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                    //                                                       .debugaccess
		.epcs_flash_controller_0_epcs_control_port_address            (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    //              epcs_flash_controller_0_epcs_control_port.address
		.epcs_flash_controller_0_epcs_control_port_write              (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),      //                                                       .write
		.epcs_flash_controller_0_epcs_control_port_read               (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),       //                                                       .read
		.epcs_flash_controller_0_epcs_control_port_readdata           (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                                                       .readdata
		.epcs_flash_controller_0_epcs_control_port_writedata          (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                                                       .writedata
		.epcs_flash_controller_0_epcs_control_port_chipselect         (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                  //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                    //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                     //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                 //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),              //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),               //                                                       .chipselect
		.LCD_RESET_N_s1_address                                       (mm_interconnect_0_lcd_reset_n_s1_address),                               //                                         LCD_RESET_N_s1.address
		.LCD_RESET_N_s1_write                                         (mm_interconnect_0_lcd_reset_n_s1_write),                                 //                                                       .write
		.LCD_RESET_N_s1_readdata                                      (mm_interconnect_0_lcd_reset_n_s1_readdata),                              //                                                       .readdata
		.LCD_RESET_N_s1_writedata                                     (mm_interconnect_0_lcd_reset_n_s1_writedata),                             //                                                       .writedata
		.LCD_RESET_N_s1_chipselect                                    (mm_interconnect_0_lcd_reset_n_s1_chipselect),                            //                                                       .chipselect
		.LT24_Controller_0_avalon_slave_0_address                     (mm_interconnect_0_lt24_controller_0_avalon_slave_0_address),             //                       LT24_Controller_0_avalon_slave_0.address
		.LT24_Controller_0_avalon_slave_0_write                       (mm_interconnect_0_lt24_controller_0_avalon_slave_0_write),               //                                                       .write
		.LT24_Controller_0_avalon_slave_0_writedata                   (mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata),           //                                                       .writedata
		.LT24_Controller_0_avalon_slave_0_chipselect                  (mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect),          //                                                       .chipselect
		.sdram_s1_address                                             (mm_interconnect_0_sdram_s1_address),                                     //                                               sdram_s1.address
		.sdram_s1_write                                               (mm_interconnect_0_sdram_s1_write),                                       //                                                       .write
		.sdram_s1_read                                                (mm_interconnect_0_sdram_s1_read),                                        //                                                       .read
		.sdram_s1_readdata                                            (mm_interconnect_0_sdram_s1_readdata),                                    //                                                       .readdata
		.sdram_s1_writedata                                           (mm_interconnect_0_sdram_s1_writedata),                                   //                                                       .writedata
		.sdram_s1_byteenable                                          (mm_interconnect_0_sdram_s1_byteenable),                                  //                                                       .byteenable
		.sdram_s1_readdatavalid                                       (mm_interconnect_0_sdram_s1_readdatavalid),                               //                                                       .readdatavalid
		.sdram_s1_waitrequest                                         (mm_interconnect_0_sdram_s1_waitrequest),                                 //                                                       .waitrequest
		.sdram_s1_chipselect                                          (mm_interconnect_0_sdram_s1_chipselect),                                  //                                                       .chipselect
		.touch_panel_busy_s1_address                                  (mm_interconnect_0_touch_panel_busy_s1_address),                          //                                    touch_panel_busy_s1.address
		.touch_panel_busy_s1_readdata                                 (mm_interconnect_0_touch_panel_busy_s1_readdata),                         //                                                       .readdata
		.touch_panel_pen_irq_n_s1_address                             (mm_interconnect_0_touch_panel_pen_irq_n_s1_address),                     //                               touch_panel_pen_irq_n_s1.address
		.touch_panel_pen_irq_n_s1_write                               (mm_interconnect_0_touch_panel_pen_irq_n_s1_write),                       //                                                       .write
		.touch_panel_pen_irq_n_s1_readdata                            (mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata),                    //                                                       .readdata
		.touch_panel_pen_irq_n_s1_writedata                           (mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata),                   //                                                       .writedata
		.touch_panel_pen_irq_n_s1_chipselect                          (mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect),                  //                                                       .chipselect
		.touch_panel_spi_spi_control_port_address                     (mm_interconnect_0_touch_panel_spi_spi_control_port_address),             //                       touch_panel_spi_spi_control_port.address
		.touch_panel_spi_spi_control_port_write                       (mm_interconnect_0_touch_panel_spi_spi_control_port_write),               //                                                       .write
		.touch_panel_spi_spi_control_port_read                        (mm_interconnect_0_touch_panel_spi_spi_control_port_read),                //                                                       .read
		.touch_panel_spi_spi_control_port_readdata                    (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),            //                                                       .readdata
		.touch_panel_spi_spi_control_port_writedata                   (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),           //                                                       .writedata
		.touch_panel_spi_spi_control_port_chipselect                  (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect)           //                                                       .chipselect
	);

	DE0_Nano_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.altpll_sys_c2_clk                                      (altpll_sys_c2_clk),                              //                                    altpll_sys_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                 // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                   //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),               //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                      //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                  //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),             //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                     //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                 //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),               //                                                 .debugaccess
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),               //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                 //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),              //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),             //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),            //                                                 .chipselect
		.led_s1_address                                         (mm_interconnect_1_led_s1_address),               //                                           led_s1.address
		.led_s1_write                                           (mm_interconnect_1_led_s1_write),                 //                                                 .write
		.led_s1_readdata                                        (mm_interconnect_1_led_s1_readdata),              //                                                 .readdata
		.led_s1_writedata                                       (mm_interconnect_1_led_s1_writedata),             //                                                 .writedata
		.led_s1_chipselect                                      (mm_interconnect_1_led_s1_chipselect),            //                                                 .chipselect
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                  //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),               //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),              //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),             //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),  //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata), //                                                 .readdata
		.timer_s1_address                                       (mm_interconnect_1_timer_s1_address),             //                                         timer_s1.address
		.timer_s1_write                                         (mm_interconnect_1_timer_s1_write),               //                                                 .write
		.timer_s1_readdata                                      (mm_interconnect_1_timer_s1_readdata),            //                                                 .readdata
		.timer_s1_writedata                                     (mm_interconnect_1_timer_s1_writedata),           //                                                 .writedata
		.timer_s1_chipselect                                    (mm_interconnect_1_timer_s1_chipselect)           //                                                 .chipselect
	);

	DE0_Nano_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_sys_c0_clk),                  //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_sys_c2_clk),                  //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_sys_c2_clk),                  //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_sys_c2_clk),                  //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                          // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_sys_c2_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (altpll_sys_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
