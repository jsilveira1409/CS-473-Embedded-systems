-- soc_system_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_tb is
end entity soc_system_tb;

architecture rtl of soc_system_tb is
	component soc_system is
		port (
			clk_clk                             : in    std_logic                     := 'X';             -- clk
			hps_0_ddr_mem_a                     : out   std_logic_vector(14 downto 0);                    -- mem_a
			hps_0_ddr_mem_ba                    : out   std_logic_vector(2 downto 0);                     -- mem_ba
			hps_0_ddr_mem_ck                    : out   std_logic;                                        -- mem_ck
			hps_0_ddr_mem_ck_n                  : out   std_logic;                                        -- mem_ck_n
			hps_0_ddr_mem_cke                   : out   std_logic;                                        -- mem_cke
			hps_0_ddr_mem_cs_n                  : out   std_logic;                                        -- mem_cs_n
			hps_0_ddr_mem_ras_n                 : out   std_logic;                                        -- mem_ras_n
			hps_0_ddr_mem_cas_n                 : out   std_logic;                                        -- mem_cas_n
			hps_0_ddr_mem_we_n                  : out   std_logic;                                        -- mem_we_n
			hps_0_ddr_mem_reset_n               : out   std_logic;                                        -- mem_reset_n
			hps_0_ddr_mem_dq                    : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			hps_0_ddr_mem_dqs                   : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			hps_0_ddr_mem_dqs_n                 : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			hps_0_ddr_mem_odt                   : out   std_logic;                                        -- mem_odt
			hps_0_ddr_mem_dm                    : out   std_logic_vector(3 downto 0);                     -- mem_dm
			hps_0_ddr_oct_rzqin                 : in    std_logic                     := 'X';             -- oct_rzqin
			hps_0_io_hps_io_emac1_inst_TX_CLK   : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_0_io_hps_io_emac1_inst_TXD0     : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_0_io_hps_io_emac1_inst_TXD1     : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_0_io_hps_io_emac1_inst_TXD2     : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_0_io_hps_io_emac1_inst_TXD3     : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_0_io_hps_io_emac1_inst_RXD0     : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_0_io_hps_io_emac1_inst_MDIO     : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_0_io_hps_io_emac1_inst_MDC      : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_0_io_hps_io_emac1_inst_RX_CTL   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_0_io_hps_io_emac1_inst_TX_CTL   : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_0_io_hps_io_emac1_inst_RX_CLK   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_0_io_hps_io_emac1_inst_RXD1     : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_0_io_hps_io_emac1_inst_RXD2     : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_0_io_hps_io_emac1_inst_RXD3     : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_0_io_hps_io_sdio_inst_CMD       : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_0_io_hps_io_sdio_inst_D0        : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_0_io_hps_io_sdio_inst_D1        : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_0_io_hps_io_sdio_inst_CLK       : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_0_io_hps_io_sdio_inst_D2        : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_0_io_hps_io_sdio_inst_D3        : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_0_io_hps_io_usb1_inst_D0        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_0_io_hps_io_usb1_inst_D1        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_0_io_hps_io_usb1_inst_D2        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_0_io_hps_io_usb1_inst_D3        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_0_io_hps_io_usb1_inst_D4        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_0_io_hps_io_usb1_inst_D5        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_0_io_hps_io_usb1_inst_D6        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_0_io_hps_io_usb1_inst_D7        : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_0_io_hps_io_usb1_inst_CLK       : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_0_io_hps_io_usb1_inst_STP       : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_0_io_hps_io_usb1_inst_DIR       : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_0_io_hps_io_usb1_inst_NXT       : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_0_io_hps_io_spim1_inst_CLK      : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_0_io_hps_io_spim1_inst_MOSI     : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_0_io_hps_io_spim1_inst_MISO     : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_0_io_hps_io_spim1_inst_SS0      : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_0_io_hps_io_uart0_inst_RX       : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_0_io_hps_io_uart0_inst_TX       : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_0_io_hps_io_i2c0_inst_SDA       : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_0_io_hps_io_i2c0_inst_SCL       : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_0_io_hps_io_i2c1_inst_SDA       : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_0_io_hps_io_i2c1_inst_SCL       : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_0_io_hps_io_gpio_inst_GPIO09    : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_0_io_hps_io_gpio_inst_GPIO35    : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_0_io_hps_io_gpio_inst_GPIO40    : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_0_io_hps_io_gpio_inst_GPIO53    : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_0_io_hps_io_gpio_inst_GPIO54    : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_0_io_hps_io_gpio_inst_GPIO61    : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			lcd_0_output_csx                    : out   std_logic;                                        -- csx
			lcd_0_output_dcx                    : out   std_logic;                                        -- dcx
			lcd_0_output_d                      : out   std_logic_vector(15 downto 0);                    -- d
			lcd_0_output_resx                   : out   std_logic;                                        -- resx
			lcd_0_output_wrx                    : out   std_logic;                                        -- wrx
			pio_leds_external_connection_export : out   std_logic_vector(7 downto 0);                     -- export
			reset_reset_n                       : in    std_logic                     := 'X'              -- reset_n
		);
	end component soc_system;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			sig_mem_a       : in    std_logic_vector(14 downto 0) := (others => 'X'); -- mem_a
			sig_mem_ba      : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- mem_ba
			sig_mem_cas_n   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cas_n
			sig_mem_ck      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_ck
			sig_mem_ck_n    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_ck_n
			sig_mem_cke     : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cke
			sig_mem_cs_n    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cs_n
			sig_mem_dm      : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dm
			sig_mem_dq      : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			sig_mem_dqs     : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			sig_mem_dqs_n   : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			sig_mem_odt     : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_odt
			sig_mem_ras_n   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_ras_n
			sig_mem_reset_n : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_reset_n
			sig_mem_we_n    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_we_n
			sig_oct_rzqin   : out   std_logic_vector(0 downto 0)                      -- oct_rzqin
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_hps_io_emac1_inst_MDC    : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_MDC
			sig_hps_io_emac1_inst_MDIO   : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_MDIO
			sig_hps_io_emac1_inst_RXD0   : out   std_logic_vector(0 downto 0);                    -- hps_io_emac1_inst_RXD0
			sig_hps_io_emac1_inst_RXD1   : out   std_logic_vector(0 downto 0);                    -- hps_io_emac1_inst_RXD1
			sig_hps_io_emac1_inst_RXD2   : out   std_logic_vector(0 downto 0);                    -- hps_io_emac1_inst_RXD2
			sig_hps_io_emac1_inst_RXD3   : out   std_logic_vector(0 downto 0);                    -- hps_io_emac1_inst_RXD3
			sig_hps_io_emac1_inst_RX_CLK : out   std_logic_vector(0 downto 0);                    -- hps_io_emac1_inst_RX_CLK
			sig_hps_io_emac1_inst_RX_CTL : out   std_logic_vector(0 downto 0);                    -- hps_io_emac1_inst_RX_CTL
			sig_hps_io_emac1_inst_TXD0   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_TXD0
			sig_hps_io_emac1_inst_TXD1   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_TXD1
			sig_hps_io_emac1_inst_TXD2   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_TXD2
			sig_hps_io_emac1_inst_TXD3   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_TXD3
			sig_hps_io_emac1_inst_TX_CLK : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_TX_CLK
			sig_hps_io_emac1_inst_TX_CTL : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_emac1_inst_TX_CTL
			sig_hps_io_gpio_inst_GPIO09  : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_gpio_inst_GPIO09
			sig_hps_io_gpio_inst_GPIO35  : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_gpio_inst_GPIO35
			sig_hps_io_gpio_inst_GPIO40  : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_gpio_inst_GPIO40
			sig_hps_io_gpio_inst_GPIO53  : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_gpio_inst_GPIO53
			sig_hps_io_gpio_inst_GPIO54  : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_gpio_inst_GPIO54
			sig_hps_io_gpio_inst_GPIO61  : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_gpio_inst_GPIO61
			sig_hps_io_i2c0_inst_SCL     : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_i2c0_inst_SCL
			sig_hps_io_i2c0_inst_SDA     : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_i2c0_inst_SDA
			sig_hps_io_i2c1_inst_SCL     : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_i2c1_inst_SCL
			sig_hps_io_i2c1_inst_SDA     : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_i2c1_inst_SDA
			sig_hps_io_sdio_inst_CLK     : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_sdio_inst_CLK
			sig_hps_io_sdio_inst_CMD     : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_sdio_inst_CMD
			sig_hps_io_sdio_inst_D0      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_sdio_inst_D0
			sig_hps_io_sdio_inst_D1      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_sdio_inst_D1
			sig_hps_io_sdio_inst_D2      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_sdio_inst_D2
			sig_hps_io_sdio_inst_D3      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_sdio_inst_D3
			sig_hps_io_spim1_inst_CLK    : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_spim1_inst_CLK
			sig_hps_io_spim1_inst_MISO   : out   std_logic_vector(0 downto 0);                    -- hps_io_spim1_inst_MISO
			sig_hps_io_spim1_inst_MOSI   : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_spim1_inst_MOSI
			sig_hps_io_spim1_inst_SS0    : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_spim1_inst_SS0
			sig_hps_io_uart0_inst_RX     : out   std_logic_vector(0 downto 0);                    -- hps_io_uart0_inst_RX
			sig_hps_io_uart0_inst_TX     : in    std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_uart0_inst_TX
			sig_hps_io_usb1_inst_CLK     : out   std_logic_vector(0 downto 0);                    -- hps_io_usb1_inst_CLK
			sig_hps_io_usb1_inst_D0      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D0
			sig_hps_io_usb1_inst_D1      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D1
			sig_hps_io_usb1_inst_D2      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D2
			sig_hps_io_usb1_inst_D3      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D3
			sig_hps_io_usb1_inst_D4      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D4
			sig_hps_io_usb1_inst_D5      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D5
			sig_hps_io_usb1_inst_D6      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D6
			sig_hps_io_usb1_inst_D7      : inout std_logic_vector(0 downto 0) := (others => 'X'); -- hps_io_usb1_inst_D7
			sig_hps_io_usb1_inst_DIR     : out   std_logic_vector(0 downto 0);                    -- hps_io_usb1_inst_DIR
			sig_hps_io_usb1_inst_NXT     : out   std_logic_vector(0 downto 0);                    -- hps_io_usb1_inst_NXT
			sig_hps_io_usb1_inst_STP     : in    std_logic_vector(0 downto 0) := (others => 'X')  -- hps_io_usb1_inst_STP
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk      : in std_logic                     := 'X';             -- clk
			reset    : in std_logic                     := 'X';             -- reset
			sig_csx  : in std_logic_vector(0 downto 0)  := (others => 'X'); -- csx
			sig_d    : in std_logic_vector(15 downto 0) := (others => 'X'); -- d
			sig_dcx  : in std_logic_vector(0 downto 0)  := (others => 'X'); -- dcx
			sig_resx : in std_logic_vector(0 downto 0)  := (others => 'X'); -- resx
			sig_wrx  : in std_logic_vector(0 downto 0)  := (others => 'X')  -- wrx
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			sig_export : in std_logic_vector(7 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0004;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal soc_system_inst_clk_bfm_clk_clk                               : std_logic;                     -- soc_system_inst_clk_bfm:clk -> [soc_system_inst:clk_clk, soc_system_inst_lcd_0_output_bfm:clk, soc_system_inst_reset_bfm:clk]
	signal soc_system_inst_hps_0_ddr_bfm_conduit_oct_rzqin               : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_ddr_bfm:sig_oct_rzqin -> soc_system_inst:hps_0_ddr_oct_rzqin
	signal soc_system_inst_hps_0_ddr_mem_cas_n                           : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_cas_n -> soc_system_inst_hps_0_ddr_bfm:sig_mem_cas_n
	signal soc_system_inst_hps_0_ddr_mem_reset_n                         : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_reset_n -> soc_system_inst_hps_0_ddr_bfm:sig_mem_reset_n
	signal soc_system_inst_hps_0_ddr_mem_ba                              : std_logic_vector(2 downto 0);  -- soc_system_inst:hps_0_ddr_mem_ba -> soc_system_inst_hps_0_ddr_bfm:sig_mem_ba
	signal soc_system_inst_hps_0_ddr_mem_we_n                            : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_we_n -> soc_system_inst_hps_0_ddr_bfm:sig_mem_we_n
	signal soc_system_inst_hps_0_ddr_mem_ck                              : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_ck -> soc_system_inst_hps_0_ddr_bfm:sig_mem_ck
	signal soc_system_inst_hps_0_ddr_mem_dm                              : std_logic_vector(3 downto 0);  -- soc_system_inst:hps_0_ddr_mem_dm -> soc_system_inst_hps_0_ddr_bfm:sig_mem_dm
	signal soc_system_inst_hps_0_ddr_mem_dqs                             : std_logic_vector(3 downto 0);  -- [] -> [soc_system_inst:hps_0_ddr_mem_dqs, soc_system_inst_hps_0_ddr_bfm:sig_mem_dqs]
	signal soc_system_inst_hps_0_ddr_mem_dq                              : std_logic_vector(31 downto 0); -- [] -> [soc_system_inst:hps_0_ddr_mem_dq, soc_system_inst_hps_0_ddr_bfm:sig_mem_dq]
	signal soc_system_inst_hps_0_ddr_mem_cs_n                            : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_cs_n -> soc_system_inst_hps_0_ddr_bfm:sig_mem_cs_n
	signal soc_system_inst_hps_0_ddr_mem_a                               : std_logic_vector(14 downto 0); -- soc_system_inst:hps_0_ddr_mem_a -> soc_system_inst_hps_0_ddr_bfm:sig_mem_a
	signal soc_system_inst_hps_0_ddr_mem_dqs_n                           : std_logic_vector(3 downto 0);  -- [] -> [soc_system_inst:hps_0_ddr_mem_dqs_n, soc_system_inst_hps_0_ddr_bfm:sig_mem_dqs_n]
	signal soc_system_inst_hps_0_ddr_mem_odt                             : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_odt -> soc_system_inst_hps_0_ddr_bfm:sig_mem_odt
	signal soc_system_inst_hps_0_ddr_mem_ras_n                           : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_ras_n -> soc_system_inst_hps_0_ddr_bfm:sig_mem_ras_n
	signal soc_system_inst_hps_0_ddr_mem_ck_n                            : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_ck_n -> soc_system_inst_hps_0_ddr_bfm:sig_mem_ck_n
	signal soc_system_inst_hps_0_ddr_mem_cke                             : std_logic;                     -- soc_system_inst:hps_0_ddr_mem_cke -> soc_system_inst_hps_0_ddr_bfm:sig_mem_cke
	signal soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio35              : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_gpio_inst_GPIO35, soc_system_inst_hps_0_io_bfm:sig_hps_io_gpio_inst_GPIO35]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_spim1_inst_miso   : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_spim1_inst_MISO -> soc_system_inst:hps_0_io_hps_io_spim1_inst_MISO
	signal soc_system_inst_hps_0_io_hps_io_spim1_inst_mosi               : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_spim1_inst_MOSI -> soc_system_inst_hps_0_io_bfm:sig_hps_io_spim1_inst_MOSI
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_mdio               : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_emac1_inst_MDIO, soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_MDIO]
	signal soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio54              : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_gpio_inst_GPIO54, soc_system_inst_hps_0_io_bfm:sig_hps_io_gpio_inst_GPIO54]
	signal soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio53              : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_gpio_inst_GPIO53, soc_system_inst_hps_0_io_bfm:sig_hps_io_gpio_inst_GPIO53]
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_tx_clk             : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_TX_CLK -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_TX_CLK
	signal soc_system_inst_hps_0_io_hps_io_i2c0_inst_scl                 : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_i2c0_inst_SCL, soc_system_inst_hps_0_io_bfm:sig_hps_io_i2c0_inst_SCL]
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_stp                 : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_usb1_inst_STP -> soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_STP
	signal soc_system_inst_hps_0_io_hps_io_sdio_inst_d3                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_sdio_inst_D3, soc_system_inst_hps_0_io_bfm:sig_hps_io_sdio_inst_D3]
	signal soc_system_inst_hps_0_io_hps_io_sdio_inst_d2                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_sdio_inst_D2, soc_system_inst_hps_0_io_bfm:sig_hps_io_sdio_inst_D2]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd3   : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_RXD3 -> soc_system_inst:hps_0_io_hps_io_emac1_inst_RXD3
	signal soc_system_inst_hps_0_io_hps_io_sdio_inst_clk                 : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_sdio_inst_CLK -> soc_system_inst_hps_0_io_bfm:sig_hps_io_sdio_inst_CLK
	signal soc_system_inst_hps_0_io_hps_io_sdio_inst_d1                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_sdio_inst_D1, soc_system_inst_hps_0_io_bfm:sig_hps_io_sdio_inst_D1]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd2   : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_RXD2 -> soc_system_inst:hps_0_io_hps_io_emac1_inst_RXD2
	signal soc_system_inst_hps_0_io_hps_io_sdio_inst_d0                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_sdio_inst_D0, soc_system_inst_hps_0_io_bfm:sig_hps_io_sdio_inst_D0]
	signal soc_system_inst_hps_0_io_hps_io_spim1_inst_clk                : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_spim1_inst_CLK -> soc_system_inst_hps_0_io_bfm:sig_hps_io_spim1_inst_CLK
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_txd2               : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_TXD2 -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_TXD2
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_txd3               : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_TXD3 -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_TXD3
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd1   : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_RXD1 -> soc_system_inst:hps_0_io_hps_io_emac1_inst_RXD1
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_txd0               : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_TXD0 -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_TXD0
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd0   : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_RXD0 -> soc_system_inst:hps_0_io_hps_io_emac1_inst_RXD0
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_txd1               : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_TXD1 -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_TXD1
	signal soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio09              : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_gpio_inst_GPIO09, soc_system_inst_hps_0_io_bfm:sig_hps_io_gpio_inst_GPIO09]
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_mdc                : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_MDC -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_MDC
	signal soc_system_inst_hps_0_io_hps_io_i2c0_inst_sda                 : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_i2c0_inst_SDA, soc_system_inst_hps_0_io_bfm:sig_hps_io_i2c0_inst_SDA]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rx_clk : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_RX_CLK -> soc_system_inst:hps_0_io_hps_io_emac1_inst_RX_CLK
	signal soc_system_inst_hps_0_io_hps_io_sdio_inst_cmd                 : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_sdio_inst_CMD, soc_system_inst_hps_0_io_bfm:sig_hps_io_sdio_inst_CMD]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_dir     : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_DIR -> soc_system_inst:hps_0_io_hps_io_usb1_inst_DIR
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rx_ctl : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_RX_CTL -> soc_system_inst:hps_0_io_hps_io_emac1_inst_RX_CTL
	signal soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio40              : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_gpio_inst_GPIO40, soc_system_inst_hps_0_io_bfm:sig_hps_io_gpio_inst_GPIO40]
	signal soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio61              : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_gpio_inst_GPIO61, soc_system_inst_hps_0_io_bfm:sig_hps_io_gpio_inst_GPIO61]
	signal soc_system_inst_hps_0_io_hps_io_i2c1_inst_scl                 : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_i2c1_inst_SCL, soc_system_inst_hps_0_io_bfm:sig_hps_io_i2c1_inst_SCL]
	signal soc_system_inst_hps_0_io_hps_io_i2c1_inst_sda                 : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_i2c1_inst_SDA, soc_system_inst_hps_0_io_bfm:sig_hps_io_i2c1_inst_SDA]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_clk     : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_CLK -> soc_system_inst:hps_0_io_hps_io_usb1_inst_CLK
	signal soc_system_inst_hps_0_io_hps_io_uart0_inst_tx                 : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_uart0_inst_TX -> soc_system_inst_hps_0_io_bfm:sig_hps_io_uart0_inst_TX
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d4                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D4, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D4]
	signal soc_system_inst_hps_0_io_hps_io_emac1_inst_tx_ctl             : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_emac1_inst_TX_CTL -> soc_system_inst_hps_0_io_bfm:sig_hps_io_emac1_inst_TX_CTL
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d5                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D5, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D5]
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d6                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D6, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D6]
	signal soc_system_inst_hps_0_io_hps_io_spim1_inst_ss0                : std_logic;                     -- soc_system_inst:hps_0_io_hps_io_spim1_inst_SS0 -> soc_system_inst_hps_0_io_bfm:sig_hps_io_spim1_inst_SS0
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d7                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D7, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D7]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_nxt     : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_NXT -> soc_system_inst:hps_0_io_hps_io_usb1_inst_NXT
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d0                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D0, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D0]
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d1                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D1, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D1]
	signal soc_system_inst_hps_0_io_bfm_conduit_hps_io_uart0_inst_rx     : std_logic_vector(0 downto 0);  -- soc_system_inst_hps_0_io_bfm:sig_hps_io_uart0_inst_RX -> soc_system_inst:hps_0_io_hps_io_uart0_inst_RX
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d2                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D2, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D2]
	signal soc_system_inst_hps_0_io_hps_io_usb1_inst_d3                  : std_logic;                     -- [] -> [soc_system_inst:hps_0_io_hps_io_usb1_inst_D3, soc_system_inst_hps_0_io_bfm:sig_hps_io_usb1_inst_D3]
	signal soc_system_inst_lcd_0_output_d                                : std_logic_vector(15 downto 0); -- soc_system_inst:lcd_0_output_d -> soc_system_inst_lcd_0_output_bfm:sig_d
	signal soc_system_inst_lcd_0_output_dcx                              : std_logic;                     -- soc_system_inst:lcd_0_output_dcx -> soc_system_inst_lcd_0_output_bfm:sig_dcx
	signal soc_system_inst_lcd_0_output_csx                              : std_logic;                     -- soc_system_inst:lcd_0_output_csx -> soc_system_inst_lcd_0_output_bfm:sig_csx
	signal soc_system_inst_lcd_0_output_wrx                              : std_logic;                     -- soc_system_inst:lcd_0_output_wrx -> soc_system_inst_lcd_0_output_bfm:sig_wrx
	signal soc_system_inst_lcd_0_output_resx                             : std_logic;                     -- soc_system_inst:lcd_0_output_resx -> soc_system_inst_lcd_0_output_bfm:sig_resx
	signal soc_system_inst_pio_leds_external_connection_export           : std_logic_vector(7 downto 0);  -- soc_system_inst:pio_leds_external_connection_export -> soc_system_inst_pio_leds_external_connection_bfm:sig_export
	signal soc_system_inst_reset_bfm_reset_reset                         : std_logic;                     -- soc_system_inst_reset_bfm:reset -> [soc_system_inst:reset_reset_n, soc_system_inst_reset_bfm_reset_reset:in]
	signal soc_system_inst_reset_bfm_reset_reset_ports_inv               : std_logic;                     -- soc_system_inst_reset_bfm_reset_reset:inv -> soc_system_inst_lcd_0_output_bfm:reset

begin

	soc_system_inst : component soc_system
		port map (
			clk_clk                             => soc_system_inst_clk_bfm_clk_clk,                                  --                          clk.clk
			hps_0_ddr_mem_a                     => soc_system_inst_hps_0_ddr_mem_a,                                  --                    hps_0_ddr.mem_a
			hps_0_ddr_mem_ba                    => soc_system_inst_hps_0_ddr_mem_ba,                                 --                             .mem_ba
			hps_0_ddr_mem_ck                    => soc_system_inst_hps_0_ddr_mem_ck,                                 --                             .mem_ck
			hps_0_ddr_mem_ck_n                  => soc_system_inst_hps_0_ddr_mem_ck_n,                               --                             .mem_ck_n
			hps_0_ddr_mem_cke                   => soc_system_inst_hps_0_ddr_mem_cke,                                --                             .mem_cke
			hps_0_ddr_mem_cs_n                  => soc_system_inst_hps_0_ddr_mem_cs_n,                               --                             .mem_cs_n
			hps_0_ddr_mem_ras_n                 => soc_system_inst_hps_0_ddr_mem_ras_n,                              --                             .mem_ras_n
			hps_0_ddr_mem_cas_n                 => soc_system_inst_hps_0_ddr_mem_cas_n,                              --                             .mem_cas_n
			hps_0_ddr_mem_we_n                  => soc_system_inst_hps_0_ddr_mem_we_n,                               --                             .mem_we_n
			hps_0_ddr_mem_reset_n               => soc_system_inst_hps_0_ddr_mem_reset_n,                            --                             .mem_reset_n
			hps_0_ddr_mem_dq                    => soc_system_inst_hps_0_ddr_mem_dq,                                 --                             .mem_dq
			hps_0_ddr_mem_dqs                   => soc_system_inst_hps_0_ddr_mem_dqs,                                --                             .mem_dqs
			hps_0_ddr_mem_dqs_n                 => soc_system_inst_hps_0_ddr_mem_dqs_n,                              --                             .mem_dqs_n
			hps_0_ddr_mem_odt                   => soc_system_inst_hps_0_ddr_mem_odt,                                --                             .mem_odt
			hps_0_ddr_mem_dm                    => soc_system_inst_hps_0_ddr_mem_dm,                                 --                             .mem_dm
			hps_0_ddr_oct_rzqin                 => soc_system_inst_hps_0_ddr_bfm_conduit_oct_rzqin(0),               --                             .oct_rzqin
			hps_0_io_hps_io_emac1_inst_TX_CLK   => soc_system_inst_hps_0_io_hps_io_emac1_inst_tx_clk,                --                     hps_0_io.hps_io_emac1_inst_TX_CLK
			hps_0_io_hps_io_emac1_inst_TXD0     => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd0,                  --                             .hps_io_emac1_inst_TXD0
			hps_0_io_hps_io_emac1_inst_TXD1     => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd1,                  --                             .hps_io_emac1_inst_TXD1
			hps_0_io_hps_io_emac1_inst_TXD2     => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd2,                  --                             .hps_io_emac1_inst_TXD2
			hps_0_io_hps_io_emac1_inst_TXD3     => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd3,                  --                             .hps_io_emac1_inst_TXD3
			hps_0_io_hps_io_emac1_inst_RXD0     => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd0(0),   --                             .hps_io_emac1_inst_RXD0
			hps_0_io_hps_io_emac1_inst_MDIO     => soc_system_inst_hps_0_io_hps_io_emac1_inst_mdio,                  --                             .hps_io_emac1_inst_MDIO
			hps_0_io_hps_io_emac1_inst_MDC      => soc_system_inst_hps_0_io_hps_io_emac1_inst_mdc,                   --                             .hps_io_emac1_inst_MDC
			hps_0_io_hps_io_emac1_inst_RX_CTL   => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rx_ctl(0), --                             .hps_io_emac1_inst_RX_CTL
			hps_0_io_hps_io_emac1_inst_TX_CTL   => soc_system_inst_hps_0_io_hps_io_emac1_inst_tx_ctl,                --                             .hps_io_emac1_inst_TX_CTL
			hps_0_io_hps_io_emac1_inst_RX_CLK   => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rx_clk(0), --                             .hps_io_emac1_inst_RX_CLK
			hps_0_io_hps_io_emac1_inst_RXD1     => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd1(0),   --                             .hps_io_emac1_inst_RXD1
			hps_0_io_hps_io_emac1_inst_RXD2     => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd2(0),   --                             .hps_io_emac1_inst_RXD2
			hps_0_io_hps_io_emac1_inst_RXD3     => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd3(0),   --                             .hps_io_emac1_inst_RXD3
			hps_0_io_hps_io_sdio_inst_CMD       => soc_system_inst_hps_0_io_hps_io_sdio_inst_cmd,                    --                             .hps_io_sdio_inst_CMD
			hps_0_io_hps_io_sdio_inst_D0        => soc_system_inst_hps_0_io_hps_io_sdio_inst_d0,                     --                             .hps_io_sdio_inst_D0
			hps_0_io_hps_io_sdio_inst_D1        => soc_system_inst_hps_0_io_hps_io_sdio_inst_d1,                     --                             .hps_io_sdio_inst_D1
			hps_0_io_hps_io_sdio_inst_CLK       => soc_system_inst_hps_0_io_hps_io_sdio_inst_clk,                    --                             .hps_io_sdio_inst_CLK
			hps_0_io_hps_io_sdio_inst_D2        => soc_system_inst_hps_0_io_hps_io_sdio_inst_d2,                     --                             .hps_io_sdio_inst_D2
			hps_0_io_hps_io_sdio_inst_D3        => soc_system_inst_hps_0_io_hps_io_sdio_inst_d3,                     --                             .hps_io_sdio_inst_D3
			hps_0_io_hps_io_usb1_inst_D0        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d0,                     --                             .hps_io_usb1_inst_D0
			hps_0_io_hps_io_usb1_inst_D1        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d1,                     --                             .hps_io_usb1_inst_D1
			hps_0_io_hps_io_usb1_inst_D2        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d2,                     --                             .hps_io_usb1_inst_D2
			hps_0_io_hps_io_usb1_inst_D3        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d3,                     --                             .hps_io_usb1_inst_D3
			hps_0_io_hps_io_usb1_inst_D4        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d4,                     --                             .hps_io_usb1_inst_D4
			hps_0_io_hps_io_usb1_inst_D5        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d5,                     --                             .hps_io_usb1_inst_D5
			hps_0_io_hps_io_usb1_inst_D6        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d6,                     --                             .hps_io_usb1_inst_D6
			hps_0_io_hps_io_usb1_inst_D7        => soc_system_inst_hps_0_io_hps_io_usb1_inst_d7,                     --                             .hps_io_usb1_inst_D7
			hps_0_io_hps_io_usb1_inst_CLK       => soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_clk(0),     --                             .hps_io_usb1_inst_CLK
			hps_0_io_hps_io_usb1_inst_STP       => soc_system_inst_hps_0_io_hps_io_usb1_inst_stp,                    --                             .hps_io_usb1_inst_STP
			hps_0_io_hps_io_usb1_inst_DIR       => soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_dir(0),     --                             .hps_io_usb1_inst_DIR
			hps_0_io_hps_io_usb1_inst_NXT       => soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_nxt(0),     --                             .hps_io_usb1_inst_NXT
			hps_0_io_hps_io_spim1_inst_CLK      => soc_system_inst_hps_0_io_hps_io_spim1_inst_clk,                   --                             .hps_io_spim1_inst_CLK
			hps_0_io_hps_io_spim1_inst_MOSI     => soc_system_inst_hps_0_io_hps_io_spim1_inst_mosi,                  --                             .hps_io_spim1_inst_MOSI
			hps_0_io_hps_io_spim1_inst_MISO     => soc_system_inst_hps_0_io_bfm_conduit_hps_io_spim1_inst_miso(0),   --                             .hps_io_spim1_inst_MISO
			hps_0_io_hps_io_spim1_inst_SS0      => soc_system_inst_hps_0_io_hps_io_spim1_inst_ss0,                   --                             .hps_io_spim1_inst_SS0
			hps_0_io_hps_io_uart0_inst_RX       => soc_system_inst_hps_0_io_bfm_conduit_hps_io_uart0_inst_rx(0),     --                             .hps_io_uart0_inst_RX
			hps_0_io_hps_io_uart0_inst_TX       => soc_system_inst_hps_0_io_hps_io_uart0_inst_tx,                    --                             .hps_io_uart0_inst_TX
			hps_0_io_hps_io_i2c0_inst_SDA       => soc_system_inst_hps_0_io_hps_io_i2c0_inst_sda,                    --                             .hps_io_i2c0_inst_SDA
			hps_0_io_hps_io_i2c0_inst_SCL       => soc_system_inst_hps_0_io_hps_io_i2c0_inst_scl,                    --                             .hps_io_i2c0_inst_SCL
			hps_0_io_hps_io_i2c1_inst_SDA       => soc_system_inst_hps_0_io_hps_io_i2c1_inst_sda,                    --                             .hps_io_i2c1_inst_SDA
			hps_0_io_hps_io_i2c1_inst_SCL       => soc_system_inst_hps_0_io_hps_io_i2c1_inst_scl,                    --                             .hps_io_i2c1_inst_SCL
			hps_0_io_hps_io_gpio_inst_GPIO09    => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio09,                 --                             .hps_io_gpio_inst_GPIO09
			hps_0_io_hps_io_gpio_inst_GPIO35    => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio35,                 --                             .hps_io_gpio_inst_GPIO35
			hps_0_io_hps_io_gpio_inst_GPIO40    => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio40,                 --                             .hps_io_gpio_inst_GPIO40
			hps_0_io_hps_io_gpio_inst_GPIO53    => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio53,                 --                             .hps_io_gpio_inst_GPIO53
			hps_0_io_hps_io_gpio_inst_GPIO54    => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio54,                 --                             .hps_io_gpio_inst_GPIO54
			hps_0_io_hps_io_gpio_inst_GPIO61    => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio61,                 --                             .hps_io_gpio_inst_GPIO61
			lcd_0_output_csx                    => soc_system_inst_lcd_0_output_csx,                                 --                 lcd_0_output.csx
			lcd_0_output_dcx                    => soc_system_inst_lcd_0_output_dcx,                                 --                             .dcx
			lcd_0_output_d                      => soc_system_inst_lcd_0_output_d,                                   --                             .d
			lcd_0_output_resx                   => soc_system_inst_lcd_0_output_resx,                                --                             .resx
			lcd_0_output_wrx                    => soc_system_inst_lcd_0_output_wrx,                                 --                             .wrx
			pio_leds_external_connection_export => soc_system_inst_pio_leds_external_connection_export,              -- pio_leds_external_connection.export
			reset_reset_n                       => soc_system_inst_reset_bfm_reset_reset                             --                        reset.reset_n
		);

	soc_system_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => soc_system_inst_clk_bfm_clk_clk  -- clk.clk
		);

	soc_system_inst_hps_0_ddr_bfm : component altera_conduit_bfm
		port map (
			sig_mem_a          => soc_system_inst_hps_0_ddr_mem_a,                 -- conduit.mem_a
			sig_mem_ba         => soc_system_inst_hps_0_ddr_mem_ba,                --        .mem_ba
			sig_mem_cas_n(0)   => soc_system_inst_hps_0_ddr_mem_cas_n,             --        .mem_cas_n
			sig_mem_ck(0)      => soc_system_inst_hps_0_ddr_mem_ck,                --        .mem_ck
			sig_mem_ck_n(0)    => soc_system_inst_hps_0_ddr_mem_ck_n,              --        .mem_ck_n
			sig_mem_cke(0)     => soc_system_inst_hps_0_ddr_mem_cke,               --        .mem_cke
			sig_mem_cs_n(0)    => soc_system_inst_hps_0_ddr_mem_cs_n,              --        .mem_cs_n
			sig_mem_dm         => soc_system_inst_hps_0_ddr_mem_dm,                --        .mem_dm
			sig_mem_dq         => soc_system_inst_hps_0_ddr_mem_dq,                --        .mem_dq
			sig_mem_dqs        => soc_system_inst_hps_0_ddr_mem_dqs,               --        .mem_dqs
			sig_mem_dqs_n      => soc_system_inst_hps_0_ddr_mem_dqs_n,             --        .mem_dqs_n
			sig_mem_odt(0)     => soc_system_inst_hps_0_ddr_mem_odt,               --        .mem_odt
			sig_mem_ras_n(0)   => soc_system_inst_hps_0_ddr_mem_ras_n,             --        .mem_ras_n
			sig_mem_reset_n(0) => soc_system_inst_hps_0_ddr_mem_reset_n,           --        .mem_reset_n
			sig_mem_we_n(0)    => soc_system_inst_hps_0_ddr_mem_we_n,              --        .mem_we_n
			sig_oct_rzqin      => soc_system_inst_hps_0_ddr_bfm_conduit_oct_rzqin  --        .oct_rzqin
		);

	soc_system_inst_hps_0_io_bfm : component altera_conduit_bfm_0002
		port map (
			sig_hps_io_emac1_inst_MDC(0)    => soc_system_inst_hps_0_io_hps_io_emac1_inst_mdc,                -- conduit.hps_io_emac1_inst_MDC
			sig_hps_io_emac1_inst_MDIO(0)   => soc_system_inst_hps_0_io_hps_io_emac1_inst_mdio,               --        .hps_io_emac1_inst_MDIO
			sig_hps_io_emac1_inst_RXD0      => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd0,   --        .hps_io_emac1_inst_RXD0
			sig_hps_io_emac1_inst_RXD1      => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd1,   --        .hps_io_emac1_inst_RXD1
			sig_hps_io_emac1_inst_RXD2      => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd2,   --        .hps_io_emac1_inst_RXD2
			sig_hps_io_emac1_inst_RXD3      => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rxd3,   --        .hps_io_emac1_inst_RXD3
			sig_hps_io_emac1_inst_RX_CLK    => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rx_clk, --        .hps_io_emac1_inst_RX_CLK
			sig_hps_io_emac1_inst_RX_CTL    => soc_system_inst_hps_0_io_bfm_conduit_hps_io_emac1_inst_rx_ctl, --        .hps_io_emac1_inst_RX_CTL
			sig_hps_io_emac1_inst_TXD0(0)   => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd0,               --        .hps_io_emac1_inst_TXD0
			sig_hps_io_emac1_inst_TXD1(0)   => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd1,               --        .hps_io_emac1_inst_TXD1
			sig_hps_io_emac1_inst_TXD2(0)   => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd2,               --        .hps_io_emac1_inst_TXD2
			sig_hps_io_emac1_inst_TXD3(0)   => soc_system_inst_hps_0_io_hps_io_emac1_inst_txd3,               --        .hps_io_emac1_inst_TXD3
			sig_hps_io_emac1_inst_TX_CLK(0) => soc_system_inst_hps_0_io_hps_io_emac1_inst_tx_clk,             --        .hps_io_emac1_inst_TX_CLK
			sig_hps_io_emac1_inst_TX_CTL(0) => soc_system_inst_hps_0_io_hps_io_emac1_inst_tx_ctl,             --        .hps_io_emac1_inst_TX_CTL
			sig_hps_io_gpio_inst_GPIO09(0)  => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio09,              --        .hps_io_gpio_inst_GPIO09
			sig_hps_io_gpio_inst_GPIO35(0)  => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio35,              --        .hps_io_gpio_inst_GPIO35
			sig_hps_io_gpio_inst_GPIO40(0)  => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio40,              --        .hps_io_gpio_inst_GPIO40
			sig_hps_io_gpio_inst_GPIO53(0)  => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio53,              --        .hps_io_gpio_inst_GPIO53
			sig_hps_io_gpio_inst_GPIO54(0)  => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio54,              --        .hps_io_gpio_inst_GPIO54
			sig_hps_io_gpio_inst_GPIO61(0)  => soc_system_inst_hps_0_io_hps_io_gpio_inst_gpio61,              --        .hps_io_gpio_inst_GPIO61
			sig_hps_io_i2c0_inst_SCL(0)     => soc_system_inst_hps_0_io_hps_io_i2c0_inst_scl,                 --        .hps_io_i2c0_inst_SCL
			sig_hps_io_i2c0_inst_SDA(0)     => soc_system_inst_hps_0_io_hps_io_i2c0_inst_sda,                 --        .hps_io_i2c0_inst_SDA
			sig_hps_io_i2c1_inst_SCL(0)     => soc_system_inst_hps_0_io_hps_io_i2c1_inst_scl,                 --        .hps_io_i2c1_inst_SCL
			sig_hps_io_i2c1_inst_SDA(0)     => soc_system_inst_hps_0_io_hps_io_i2c1_inst_sda,                 --        .hps_io_i2c1_inst_SDA
			sig_hps_io_sdio_inst_CLK(0)     => soc_system_inst_hps_0_io_hps_io_sdio_inst_clk,                 --        .hps_io_sdio_inst_CLK
			sig_hps_io_sdio_inst_CMD(0)     => soc_system_inst_hps_0_io_hps_io_sdio_inst_cmd,                 --        .hps_io_sdio_inst_CMD
			sig_hps_io_sdio_inst_D0(0)      => soc_system_inst_hps_0_io_hps_io_sdio_inst_d0,                  --        .hps_io_sdio_inst_D0
			sig_hps_io_sdio_inst_D1(0)      => soc_system_inst_hps_0_io_hps_io_sdio_inst_d1,                  --        .hps_io_sdio_inst_D1
			sig_hps_io_sdio_inst_D2(0)      => soc_system_inst_hps_0_io_hps_io_sdio_inst_d2,                  --        .hps_io_sdio_inst_D2
			sig_hps_io_sdio_inst_D3(0)      => soc_system_inst_hps_0_io_hps_io_sdio_inst_d3,                  --        .hps_io_sdio_inst_D3
			sig_hps_io_spim1_inst_CLK(0)    => soc_system_inst_hps_0_io_hps_io_spim1_inst_clk,                --        .hps_io_spim1_inst_CLK
			sig_hps_io_spim1_inst_MISO      => soc_system_inst_hps_0_io_bfm_conduit_hps_io_spim1_inst_miso,   --        .hps_io_spim1_inst_MISO
			sig_hps_io_spim1_inst_MOSI(0)   => soc_system_inst_hps_0_io_hps_io_spim1_inst_mosi,               --        .hps_io_spim1_inst_MOSI
			sig_hps_io_spim1_inst_SS0(0)    => soc_system_inst_hps_0_io_hps_io_spim1_inst_ss0,                --        .hps_io_spim1_inst_SS0
			sig_hps_io_uart0_inst_RX        => soc_system_inst_hps_0_io_bfm_conduit_hps_io_uart0_inst_rx,     --        .hps_io_uart0_inst_RX
			sig_hps_io_uart0_inst_TX(0)     => soc_system_inst_hps_0_io_hps_io_uart0_inst_tx,                 --        .hps_io_uart0_inst_TX
			sig_hps_io_usb1_inst_CLK        => soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_clk,     --        .hps_io_usb1_inst_CLK
			sig_hps_io_usb1_inst_D0(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d0,                  --        .hps_io_usb1_inst_D0
			sig_hps_io_usb1_inst_D1(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d1,                  --        .hps_io_usb1_inst_D1
			sig_hps_io_usb1_inst_D2(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d2,                  --        .hps_io_usb1_inst_D2
			sig_hps_io_usb1_inst_D3(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d3,                  --        .hps_io_usb1_inst_D3
			sig_hps_io_usb1_inst_D4(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d4,                  --        .hps_io_usb1_inst_D4
			sig_hps_io_usb1_inst_D5(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d5,                  --        .hps_io_usb1_inst_D5
			sig_hps_io_usb1_inst_D6(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d6,                  --        .hps_io_usb1_inst_D6
			sig_hps_io_usb1_inst_D7(0)      => soc_system_inst_hps_0_io_hps_io_usb1_inst_d7,                  --        .hps_io_usb1_inst_D7
			sig_hps_io_usb1_inst_DIR        => soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_dir,     --        .hps_io_usb1_inst_DIR
			sig_hps_io_usb1_inst_NXT        => soc_system_inst_hps_0_io_bfm_conduit_hps_io_usb1_inst_nxt,     --        .hps_io_usb1_inst_NXT
			sig_hps_io_usb1_inst_STP(0)     => soc_system_inst_hps_0_io_hps_io_usb1_inst_stp                  --        .hps_io_usb1_inst_STP
		);

	soc_system_inst_lcd_0_output_bfm : component altera_conduit_bfm_0003
		port map (
			clk         => soc_system_inst_clk_bfm_clk_clk,                 --     clk.clk
			reset       => soc_system_inst_reset_bfm_reset_reset_ports_inv, --   reset.reset
			sig_csx(0)  => soc_system_inst_lcd_0_output_csx,                -- conduit.csx
			sig_d       => soc_system_inst_lcd_0_output_d,                  --        .d
			sig_dcx(0)  => soc_system_inst_lcd_0_output_dcx,                --        .dcx
			sig_resx(0) => soc_system_inst_lcd_0_output_resx,               --        .resx
			sig_wrx(0)  => soc_system_inst_lcd_0_output_wrx                 --        .wrx
		);

	soc_system_inst_pio_leds_external_connection_bfm : component altera_conduit_bfm_0004
		port map (
			sig_export => soc_system_inst_pio_leds_external_connection_export  -- conduit.export
		);

	soc_system_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => soc_system_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => soc_system_inst_clk_bfm_clk_clk        --   clk.clk
		);

	soc_system_inst_reset_bfm_reset_reset_ports_inv <= not soc_system_inst_reset_bfm_reset_reset;

end architecture rtl; -- of soc_system_tb
