
module system2 (
	clk_clk);	

	input		clk_clk;
endmodule
