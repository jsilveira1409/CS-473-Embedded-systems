// lt24_qsys.v

// Generated using ACDS version 13.1 182 at 2014.06.23.08:45:01

`timescale 1 ps / 1 ps
module lt24_qsys (
		input  wire        clk_clk,                                                 //                                       clk.clk
		input  wire        reset_reset_n,                                           //                                     reset.reset_n
		output wire        lcd_reset_n_export,                                      //                               lcd_reset_n.export
		input  wire        touch_panel_pen_irq_n_external_connection_export,        // touch_panel_pen_irq_n_external_connection.export
		input  wire        touch_panel_busy_external_connection_export,             //      touch_panel_busy_external_connection.export
		input  wire        touch_panel_spi_external_MISO,                           //                  touch_panel_spi_external.MISO
		output wire        touch_panel_spi_external_MOSI,                           //                                          .MOSI
		output wire        touch_panel_spi_external_SCLK,                           //                                          .SCLK
		output wire        touch_panel_spi_external_SS_n,                           //                                          .SS_n
		input  wire [3:0]  key_external_connection_export,                          //                   key_external_connection.export
		output wire        lt24_controller_0_conduit_end_cs,                        //             lt24_controller_0_conduit_end.cs
		output wire        lt24_controller_0_conduit_end_rs,                        //                                          .rs
		output wire        lt24_controller_0_conduit_end_rd,                        //                                          .rd
		output wire        lt24_controller_0_conduit_end_wr,                        //                                          .wr
		output wire [15:0] lt24_controller_0_conduit_end_data,                      //                                          .data
		output wire        pll_qsys_locked_export,                                  //                           pll_qsys_locked.export
		inout  wire [15:0] tristate_conduit_bridge_out_sram_tcm_data_out,           //               tristate_conduit_bridge_out.sram_tcm_data_out
		output wire [18:0] tristate_conduit_bridge_out_sram_tcm_address_out,        //                                          .sram_tcm_address_out
		output wire [0:0]  tristate_conduit_bridge_out_sram_tcm_outputenable_n_out, //                                          .sram_tcm_outputenable_n_out
		output wire [0:0]  tristate_conduit_bridge_out_sram_tcm_chipselect_n_out,   //                                          .sram_tcm_chipselect_n_out
		output wire [1:0]  tristate_conduit_bridge_out_sram_tcm_byteenable_n_out,   //                                          .sram_tcm_byteenable_n_out
		output wire [0:0]  tristate_conduit_bridge_out_sram_tcm_write_n_out         //                                          .sram_tcm_write_n_out
	);

	wire         pll_qsys_outclk0_clk;                                                 // pll_qsys:outclk_0 -> [LCD_RESET_N:clk, LT24_Controller_0:clk, irq_mapper:clk, jtag_uart:clk, key:clk, mm_interconnect_0:pll_qsys_outclk0_clk, nios2_qsys:clk, rst_controller:clk, rst_controller_001:clk, sram:clk_clk, sysid_qsys:clock, timer:clk, touch_panel_busy:clk, touch_panel_pen_irq_n:clk, touch_panel_spi:clk, tristate_conduit_bridge:clk, tristate_conduit_pin_sharer_sram:clk_clk]
	wire         sram_tcm_chipselect_n_out;                                            // sram:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_sram:tcs0_chipselect_n_out
	wire         sram_tcm_grant;                                                       // tristate_conduit_pin_sharer_sram:tcs0_grant -> sram:tcm_grant
	wire         sram_tcm_data_outen;                                                  // sram:tcm_data_outen -> tristate_conduit_pin_sharer_sram:tcs0_data_outen
	wire         sram_tcm_outputenable_n_out;                                          // sram:tcm_outputenable_n_out -> tristate_conduit_pin_sharer_sram:tcs0_outputenable_n_out
	wire         sram_tcm_request;                                                     // sram:tcm_request -> tristate_conduit_pin_sharer_sram:tcs0_request
	wire  [15:0] sram_tcm_data_out;                                                    // sram:tcm_data_out -> tristate_conduit_pin_sharer_sram:tcs0_data_out
	wire         sram_tcm_write_n_out;                                                 // sram:tcm_write_n_out -> tristate_conduit_pin_sharer_sram:tcs0_write_n_out
	wire  [18:0] sram_tcm_address_out;                                                 // sram:tcm_address_out -> tristate_conduit_pin_sharer_sram:tcs0_address_out
	wire  [15:0] sram_tcm_data_in;                                                     // tristate_conduit_pin_sharer_sram:tcs0_data_in -> sram:tcm_data_in
	wire   [1:0] sram_tcm_byteenable_n_out;                                            // sram:tcm_byteenable_n_out -> tristate_conduit_pin_sharer_sram:tcs0_byteenable_n_out
	wire   [0:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_write_n_out_out;        // tristate_conduit_pin_sharer_sram:sram_tcm_write_n_out -> tristate_conduit_bridge:tcs_sram_tcm_write_n_out
	wire  [18:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_address_out_out;        // tristate_conduit_pin_sharer_sram:sram_tcm_address_out -> tristate_conduit_bridge:tcs_sram_tcm_address_out
	wire         tristate_conduit_pin_sharer_sram_tcm_grant;                           // tristate_conduit_bridge:grant -> tristate_conduit_pin_sharer_sram:grant
	wire         tristate_conduit_pin_sharer_sram_tcm_request;                         // tristate_conduit_pin_sharer_sram:request -> tristate_conduit_bridge:request
	wire   [1:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_byteenable_n_out_out;   // tristate_conduit_pin_sharer_sram:sram_tcm_byteenable_n_out -> tristate_conduit_bridge:tcs_sram_tcm_byteenable_n_out
	wire   [0:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_outputenable_n_out_out; // tristate_conduit_pin_sharer_sram:sram_tcm_outputenable_n_out -> tristate_conduit_bridge:tcs_sram_tcm_outputenable_n_out
	wire         tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_outen;         // tristate_conduit_pin_sharer_sram:sram_tcm_data_outen -> tristate_conduit_bridge:tcs_sram_tcm_data_outen
	wire  [15:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_in;            // tristate_conduit_bridge:tcs_sram_tcm_data_in -> tristate_conduit_pin_sharer_sram:sram_tcm_data_in
	wire  [15:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_out;           // tristate_conduit_pin_sharer_sram:sram_tcm_data_out -> tristate_conduit_bridge:tcs_sram_tcm_data_out
	wire   [0:0] tristate_conduit_pin_sharer_sram_tcm_sram_tcm_chipselect_n_out_out;   // tristate_conduit_pin_sharer_sram:sram_tcm_chipselect_n_out -> tristate_conduit_bridge:tcs_sram_tcm_chipselect_n_out
	wire         nios2_qsys_jtag_debug_module_reset_reset;                             // nios2_qsys:jtag_debug_module_resetrequest -> [mm_interconnect_0:sram_reset_reset_bridge_in_reset_reset, rst_controller:reset_in1, sram:reset_reset]
	wire  [31:0] mm_interconnect_0_lcd_reset_n_s1_writedata;                           // mm_interconnect_0:LCD_RESET_N_s1_writedata -> LCD_RESET_N:writedata
	wire   [1:0] mm_interconnect_0_lcd_reset_n_s1_address;                             // mm_interconnect_0:LCD_RESET_N_s1_address -> LCD_RESET_N:address
	wire         mm_interconnect_0_lcd_reset_n_s1_chipselect;                          // mm_interconnect_0:LCD_RESET_N_s1_chipselect -> LCD_RESET_N:chipselect
	wire         mm_interconnect_0_lcd_reset_n_s1_write;                               // mm_interconnect_0:LCD_RESET_N_s1_write -> LCD_RESET_N:write_n
	wire  [31:0] mm_interconnect_0_lcd_reset_n_s1_readdata;                            // LCD_RESET_N:readdata -> mm_interconnect_0:LCD_RESET_N_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_panel_busy_s1_address;                        // mm_interconnect_0:touch_panel_busy_s1_address -> touch_panel_busy:address
	wire  [31:0] mm_interconnect_0_touch_panel_busy_s1_readdata;                       // touch_panel_busy:readdata -> mm_interconnect_0:touch_panel_busy_s1_readdata
	wire  [31:0] mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata;         // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_writedata -> LT24_Controller_0:s_writedata
	wire   [0:0] mm_interconnect_0_lt24_controller_0_avalon_slave_0_address;           // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_address -> LT24_Controller_0:s_address
	wire         mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect;        // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_chipselect -> LT24_Controller_0:s_chipselect_n
	wire         mm_interconnect_0_lt24_controller_0_avalon_slave_0_write;             // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_write -> LT24_Controller_0:s_write_n
	wire         nios2_qsys_data_master_waitrequest;                                   // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                                     // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [20:0] nios2_qsys_data_master_address;                                       // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire         nios2_qsys_data_master_write;                                         // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire         nios2_qsys_data_master_read;                                          // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire  [31:0] nios2_qsys_data_master_readdata;                                      // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                                   // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                                 // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                                    // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest;           // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;             // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;               // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_write;                 // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_read;                  // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;              // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess;           // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;            // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire         mm_interconnect_0_sram_uas_waitrequest;                               // sram:uas_waitrequest -> mm_interconnect_0:sram_uas_waitrequest
	wire   [1:0] mm_interconnect_0_sram_uas_burstcount;                                // mm_interconnect_0:sram_uas_burstcount -> sram:uas_burstcount
	wire  [15:0] mm_interconnect_0_sram_uas_writedata;                                 // mm_interconnect_0:sram_uas_writedata -> sram:uas_writedata
	wire  [18:0] mm_interconnect_0_sram_uas_address;                                   // mm_interconnect_0:sram_uas_address -> sram:uas_address
	wire         mm_interconnect_0_sram_uas_lock;                                      // mm_interconnect_0:sram_uas_lock -> sram:uas_lock
	wire         mm_interconnect_0_sram_uas_write;                                     // mm_interconnect_0:sram_uas_write -> sram:uas_write
	wire         mm_interconnect_0_sram_uas_read;                                      // mm_interconnect_0:sram_uas_read -> sram:uas_read
	wire  [15:0] mm_interconnect_0_sram_uas_readdata;                                  // sram:uas_readdata -> mm_interconnect_0:sram_uas_readdata
	wire         mm_interconnect_0_sram_uas_debugaccess;                               // mm_interconnect_0:sram_uas_debugaccess -> sram:uas_debugaccess
	wire         mm_interconnect_0_sram_uas_readdatavalid;                             // sram:uas_readdatavalid -> mm_interconnect_0:sram_uas_readdatavalid
	wire   [1:0] mm_interconnect_0_sram_uas_byteenable;                                // mm_interconnect_0:sram_uas_byteenable -> sram:uas_byteenable
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                   // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                  // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire  [31:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata;                 // mm_interconnect_0:touch_panel_pen_irq_n_s1_writedata -> touch_panel_pen_irq_n:writedata
	wire   [1:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_address;                   // mm_interconnect_0:touch_panel_pen_irq_n_s1_address -> touch_panel_pen_irq_n:address
	wire         mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect;                // mm_interconnect_0:touch_panel_pen_irq_n_s1_chipselect -> touch_panel_pen_irq_n:chipselect
	wire         mm_interconnect_0_touch_panel_pen_irq_n_s1_write;                     // mm_interconnect_0:touch_panel_pen_irq_n_s1_write -> touch_panel_pen_irq_n:write_n
	wire  [31:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata;                  // touch_panel_pen_irq_n:readdata -> mm_interconnect_0:touch_panel_pen_irq_n_s1_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                            // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [20:0] nios2_qsys_instruction_master_address;                                // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                                   // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                               // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                          // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                     // mm_interconnect_0:key_s1_address -> key:address
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                    // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                 // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                   // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                                // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                                     // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                  // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_writedata;         // mm_interconnect_0:touch_panel_spi_spi_control_port_writedata -> touch_panel_spi:data_from_cpu
	wire   [2:0] mm_interconnect_0_touch_panel_spi_spi_control_port_address;           // mm_interconnect_0:touch_panel_spi_spi_control_port_address -> touch_panel_spi:mem_addr
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect;        // mm_interconnect_0:touch_panel_spi_spi_control_port_chipselect -> touch_panel_spi:spi_select
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_write;             // mm_interconnect_0:touch_panel_spi_spi_control_port_write -> touch_panel_spi:write_n
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_read;              // mm_interconnect_0:touch_panel_spi_spi_control_port_read -> touch_panel_spi:read_n
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_readdata;          // touch_panel_spi:data_to_cpu -> mm_interconnect_0:touch_panel_spi_spi_control_port_readdata
	wire         irq_mapper_receiver0_irq;                                             // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                             // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                             // touch_panel_spi:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                             // touch_panel_pen_irq_n:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                                 // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n, rst_translator:in_reset, tristate_conduit_bridge:reset, tristate_conduit_pin_sharer_sram:reset_reset]
	wire         rst_controller_reset_out_reset_req;                                   // rst_controller:reset_req -> [nios2_qsys:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [LCD_RESET_N:reset_n, LT24_Controller_0:reset_n, jtag_uart:rst_n, key:reset_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, sysid_qsys:reset_n, timer:reset_n, touch_panel_busy:reset_n, touch_panel_pen_irq_n:reset_n, touch_panel_spi:reset_n]
	wire         rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> pll_qsys:rst

	lt24_qsys_nios2_qsys nios2_qsys (
		.clk                                   (pll_qsys_outclk0_clk),                                       //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	lt24_qsys_jtag_uart jtag_uart (
		.clk            (pll_qsys_outclk0_clk),                                      //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	lt24_qsys_LCD_RESET_N lcd_reset_n (
		.clk        (pll_qsys_outclk0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_lcd_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_reset_n_s1_readdata),   //                    .readdata
		.out_port   (lcd_reset_n_export)                           // external_connection.export
	);

	lt24_qsys_timer timer (
		.clk        (pll_qsys_outclk0_clk),                  //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	lt24_qsys_touch_panel_spi touch_panel_spi (
		.clk           (pll_qsys_outclk0_clk),                                          //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                           //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_touch_panel_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_touch_panel_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                      //              irq.irq
		.MISO          (touch_panel_spi_external_MISO),                                 //         external.export
		.MOSI          (touch_panel_spi_external_MOSI),                                 //                 .export
		.SCLK          (touch_panel_spi_external_SCLK),                                 //                 .export
		.SS_n          (touch_panel_spi_external_SS_n)                                  //                 .export
	);

	lt24_qsys_touch_panel_pen_irq_n touch_panel_pen_irq_n (
		.clk        (pll_qsys_outclk0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_touch_panel_pen_irq_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_panel_pen_irq_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata),   //                    .readdata
		.in_port    (touch_panel_pen_irq_n_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                               //                 irq.irq
	);

	lt24_qsys_touch_panel_busy touch_panel_busy (
		.clk      (pll_qsys_outclk0_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_touch_panel_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touch_panel_busy_s1_readdata), //                    .readdata
		.in_port  (touch_panel_busy_external_connection_export)     // external_connection.export
	);

	lt24_qsys_key key (
		.clk      (pll_qsys_outclk0_clk),                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	LT24_Controller lt24_controller_0 (
		.clk            (pll_qsys_outclk0_clk),                                           //          clock.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                            //          reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect_n
		.s_write_n      (~mm_interconnect_0_lt24_controller_0_avalon_slave_0_write),      //               .write_n
		.s_writedata    (mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata),   //               .writedata
		.s_address      (mm_interconnect_0_lt24_controller_0_avalon_slave_0_address),     //               .address
		.lt24_cs        (lt24_controller_0_conduit_end_cs),                               //    conduit_end.export
		.lt24_rs        (lt24_controller_0_conduit_end_rs),                               //               .export
		.lt24_rd        (lt24_controller_0_conduit_end_rd),                               //               .export
		.lt24_wr        (lt24_controller_0_conduit_end_wr),                               //               .export
		.lt24_data      (lt24_controller_0_conduit_end_data)                              //               .export
	);

	lt24_qsys_sysid_qsys sysid_qsys (
		.clock    (pll_qsys_outclk0_clk),                                //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	lt24_qsys_pll_qsys pll_qsys (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_002_reset_out_reset), //   reset.reset
		.outclk_0 (pll_qsys_outclk0_clk),               // outclk0.clk
		.locked   (pll_qsys_locked_export)              //  locked.export
	);

	lt24_qsys_sram #(
		.TCM_ADDRESS_W                  (19),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (10),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (10),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram (
		.clk_clk                (pll_qsys_outclk0_clk),                     //   clk.clk
		.reset_reset            (nios2_qsys_jtag_debug_module_reset_reset), // reset.reset
		.uas_address            (mm_interconnect_0_sram_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_0_sram_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_0_sram_uas_read),          //      .read
		.uas_write              (mm_interconnect_0_sram_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_0_sram_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_0_sram_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_0_sram_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_0_sram_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_0_sram_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_0_sram_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_0_sram_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (sram_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (sram_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (sram_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request            (sram_tcm_request),                         //      .request
		.tcm_grant              (sram_tcm_grant),                           //      .grant
		.tcm_address_out        (sram_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out   (sram_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out           (sram_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (sram_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (sram_tcm_data_in)                          //      .data_in
	);

	lt24_qsys_tristate_conduit_pin_sharer_sram tristate_conduit_pin_sharer_sram (
		.clk_clk                     (pll_qsys_outclk0_clk),                                                 //   clk.clk
		.reset_reset                 (rst_controller_reset_out_reset),                                       // reset.reset
		.request                     (tristate_conduit_pin_sharer_sram_tcm_request),                         //   tcm.request
		.grant                       (tristate_conduit_pin_sharer_sram_tcm_grant),                           //      .grant
		.sram_tcm_address_out        (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_address_out_out),        //      .sram_tcm_address_out_out
		.sram_tcm_outputenable_n_out (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_outputenable_n_out_out), //      .sram_tcm_outputenable_n_out_out
		.sram_tcm_byteenable_n_out   (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_byteenable_n_out_out),   //      .sram_tcm_byteenable_n_out_out
		.sram_tcm_write_n_out        (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_write_n_out_out),        //      .sram_tcm_write_n_out_out
		.sram_tcm_data_out           (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_out),           //      .sram_tcm_data_out_out
		.sram_tcm_data_in            (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_in),            //      .sram_tcm_data_out_in
		.sram_tcm_data_outen         (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_outen),         //      .sram_tcm_data_out_outen
		.sram_tcm_chipselect_n_out   (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_chipselect_n_out_out),   //      .sram_tcm_chipselect_n_out_out
		.tcs0_request                (sram_tcm_request),                                                     //  tcs0.request
		.tcs0_grant                  (sram_tcm_grant),                                                       //      .grant
		.tcs0_address_out            (sram_tcm_address_out),                                                 //      .address_out
		.tcs0_outputenable_n_out     (sram_tcm_outputenable_n_out),                                          //      .outputenable_n_out
		.tcs0_byteenable_n_out       (sram_tcm_byteenable_n_out),                                            //      .byteenable_n_out
		.tcs0_write_n_out            (sram_tcm_write_n_out),                                                 //      .write_n_out
		.tcs0_data_out               (sram_tcm_data_out),                                                    //      .data_out
		.tcs0_data_in                (sram_tcm_data_in),                                                     //      .data_in
		.tcs0_data_outen             (sram_tcm_data_outen),                                                  //      .data_outen
		.tcs0_chipselect_n_out       (sram_tcm_chipselect_n_out)                                             //      .chipselect_n_out
	);

	lt24_qsys_tristate_conduit_bridge tristate_conduit_bridge (
		.clk                             (pll_qsys_outclk0_clk),                                                 //   clk.clk
		.reset                           (rst_controller_reset_out_reset),                                       // reset.reset
		.request                         (tristate_conduit_pin_sharer_sram_tcm_request),                         //   tcs.request
		.grant                           (tristate_conduit_pin_sharer_sram_tcm_grant),                           //      .grant
		.tcs_sram_tcm_data_out           (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_out),           //      .sram_tcm_data_out_out
		.tcs_sram_tcm_data_outen         (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_outen),         //      .sram_tcm_data_out_outen
		.tcs_sram_tcm_data_in            (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_data_out_in),            //      .sram_tcm_data_out_in
		.tcs_sram_tcm_address_out        (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_address_out_out),        //      .sram_tcm_address_out_out
		.tcs_sram_tcm_outputenable_n_out (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_outputenable_n_out_out), //      .sram_tcm_outputenable_n_out_out
		.tcs_sram_tcm_chipselect_n_out   (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_chipselect_n_out_out),   //      .sram_tcm_chipselect_n_out_out
		.tcs_sram_tcm_byteenable_n_out   (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_byteenable_n_out_out),   //      .sram_tcm_byteenable_n_out_out
		.tcs_sram_tcm_write_n_out        (tristate_conduit_pin_sharer_sram_tcm_sram_tcm_write_n_out_out),        //      .sram_tcm_write_n_out_out
		.sram_tcm_data_out               (tristate_conduit_bridge_out_sram_tcm_data_out),                        //   out.sram_tcm_data_out
		.sram_tcm_address_out            (tristate_conduit_bridge_out_sram_tcm_address_out),                     //      .sram_tcm_address_out
		.sram_tcm_outputenable_n_out     (tristate_conduit_bridge_out_sram_tcm_outputenable_n_out),              //      .sram_tcm_outputenable_n_out
		.sram_tcm_chipselect_n_out       (tristate_conduit_bridge_out_sram_tcm_chipselect_n_out),                //      .sram_tcm_chipselect_n_out
		.sram_tcm_byteenable_n_out       (tristate_conduit_bridge_out_sram_tcm_byteenable_n_out),                //      .sram_tcm_byteenable_n_out
		.sram_tcm_write_n_out            (tristate_conduit_bridge_out_sram_tcm_write_n_out)                      //      .sram_tcm_write_n_out
	);

	lt24_qsys_mm_interconnect_0 mm_interconnect_0 (
		.pll_qsys_outclk0_clk                           (pll_qsys_outclk0_clk),                                          //                         pll_qsys_outclk0.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                            //    jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.sram_reset_reset_bridge_in_reset_reset         (nios2_qsys_jtag_debug_module_reset_reset),                      //         sram_reset_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                 (nios2_qsys_data_master_address),                                //                   nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest             (nios2_qsys_data_master_waitrequest),                            //                                         .waitrequest
		.nios2_qsys_data_master_byteenable              (nios2_qsys_data_master_byteenable),                             //                                         .byteenable
		.nios2_qsys_data_master_read                    (nios2_qsys_data_master_read),                                   //                                         .read
		.nios2_qsys_data_master_readdata                (nios2_qsys_data_master_readdata),                               //                                         .readdata
		.nios2_qsys_data_master_readdatavalid           (nios2_qsys_data_master_readdatavalid),                          //                                         .readdatavalid
		.nios2_qsys_data_master_write                   (nios2_qsys_data_master_write),                                  //                                         .write
		.nios2_qsys_data_master_writedata               (nios2_qsys_data_master_writedata),                              //                                         .writedata
		.nios2_qsys_data_master_debugaccess             (nios2_qsys_data_master_debugaccess),                            //                                         .debugaccess
		.nios2_qsys_instruction_master_address          (nios2_qsys_instruction_master_address),                         //            nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest      (nios2_qsys_instruction_master_waitrequest),                     //                                         .waitrequest
		.nios2_qsys_instruction_master_read             (nios2_qsys_instruction_master_read),                            //                                         .read
		.nios2_qsys_instruction_master_readdata         (nios2_qsys_instruction_master_readdata),                        //                                         .readdata
		.nios2_qsys_instruction_master_readdatavalid    (nios2_qsys_instruction_master_readdatavalid),                   //                                         .readdatavalid
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                         .chipselect
		.key_s1_address                                 (mm_interconnect_0_key_s1_address),                              //                                   key_s1.address
		.key_s1_readdata                                (mm_interconnect_0_key_s1_readdata),                             //                                         .readdata
		.LCD_RESET_N_s1_address                         (mm_interconnect_0_lcd_reset_n_s1_address),                      //                           LCD_RESET_N_s1.address
		.LCD_RESET_N_s1_write                           (mm_interconnect_0_lcd_reset_n_s1_write),                        //                                         .write
		.LCD_RESET_N_s1_readdata                        (mm_interconnect_0_lcd_reset_n_s1_readdata),                     //                                         .readdata
		.LCD_RESET_N_s1_writedata                       (mm_interconnect_0_lcd_reset_n_s1_writedata),                    //                                         .writedata
		.LCD_RESET_N_s1_chipselect                      (mm_interconnect_0_lcd_reset_n_s1_chipselect),                   //                                         .chipselect
		.LT24_Controller_0_avalon_slave_0_address       (mm_interconnect_0_lt24_controller_0_avalon_slave_0_address),    //         LT24_Controller_0_avalon_slave_0.address
		.LT24_Controller_0_avalon_slave_0_write         (mm_interconnect_0_lt24_controller_0_avalon_slave_0_write),      //                                         .write
		.LT24_Controller_0_avalon_slave_0_writedata     (mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata),  //                                         .writedata
		.LT24_Controller_0_avalon_slave_0_chipselect    (mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect), //                                         .chipselect
		.nios2_qsys_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),        //             nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),          //                                         .write
		.nios2_qsys_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),           //                                         .read
		.nios2_qsys_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),       //                                         .readdata
		.nios2_qsys_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),      //                                         .writedata
		.nios2_qsys_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),     //                                         .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest),    //                                         .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess),    //                                         .debugaccess
		.sram_uas_address                               (mm_interconnect_0_sram_uas_address),                            //                                 sram_uas.address
		.sram_uas_write                                 (mm_interconnect_0_sram_uas_write),                              //                                         .write
		.sram_uas_read                                  (mm_interconnect_0_sram_uas_read),                               //                                         .read
		.sram_uas_readdata                              (mm_interconnect_0_sram_uas_readdata),                           //                                         .readdata
		.sram_uas_writedata                             (mm_interconnect_0_sram_uas_writedata),                          //                                         .writedata
		.sram_uas_burstcount                            (mm_interconnect_0_sram_uas_burstcount),                         //                                         .burstcount
		.sram_uas_byteenable                            (mm_interconnect_0_sram_uas_byteenable),                         //                                         .byteenable
		.sram_uas_readdatavalid                         (mm_interconnect_0_sram_uas_readdatavalid),                      //                                         .readdatavalid
		.sram_uas_waitrequest                           (mm_interconnect_0_sram_uas_waitrequest),                        //                                         .waitrequest
		.sram_uas_lock                                  (mm_interconnect_0_sram_uas_lock),                               //                                         .lock
		.sram_uas_debugaccess                           (mm_interconnect_0_sram_uas_debugaccess),                        //                                         .debugaccess
		.sysid_qsys_control_slave_address               (mm_interconnect_0_sysid_qsys_control_slave_address),            //                 sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata              (mm_interconnect_0_sysid_qsys_control_slave_readdata),           //                                         .readdata
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                            //                                 timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                              //                                         .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                           //                                         .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                          //                                         .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect),                         //                                         .chipselect
		.touch_panel_busy_s1_address                    (mm_interconnect_0_touch_panel_busy_s1_address),                 //                      touch_panel_busy_s1.address
		.touch_panel_busy_s1_readdata                   (mm_interconnect_0_touch_panel_busy_s1_readdata),                //                                         .readdata
		.touch_panel_pen_irq_n_s1_address               (mm_interconnect_0_touch_panel_pen_irq_n_s1_address),            //                 touch_panel_pen_irq_n_s1.address
		.touch_panel_pen_irq_n_s1_write                 (mm_interconnect_0_touch_panel_pen_irq_n_s1_write),              //                                         .write
		.touch_panel_pen_irq_n_s1_readdata              (mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata),           //                                         .readdata
		.touch_panel_pen_irq_n_s1_writedata             (mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata),          //                                         .writedata
		.touch_panel_pen_irq_n_s1_chipselect            (mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect),         //                                         .chipselect
		.touch_panel_spi_spi_control_port_address       (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //         touch_panel_spi_spi_control_port.address
		.touch_panel_spi_spi_control_port_write         (mm_interconnect_0_touch_panel_spi_spi_control_port_write),      //                                         .write
		.touch_panel_spi_spi_control_port_read          (mm_interconnect_0_touch_panel_spi_spi_control_port_read),       //                                         .read
		.touch_panel_spi_spi_control_port_readdata      (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                                         .readdata
		.touch_panel_spi_spi_control_port_writedata     (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  //                                         .writedata
		.touch_panel_spi_spi_control_port_chipselect    (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect)  //                                         .chipselect
	);

	lt24_qsys_irq_mapper irq_mapper (
		.clk           (pll_qsys_outclk0_clk),           //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (pll_qsys_outclk0_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_qsys_outclk0_clk),               //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
