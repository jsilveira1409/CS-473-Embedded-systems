
module system (
	clk_clk,
	daisyport_0_conduit_end_writeresponsevalid_n,
	reset_reset_n);	

	input		clk_clk;
	output		daisyport_0_conduit_end_writeresponsevalid_n;
	input		reset_reset_n;
endmodule
