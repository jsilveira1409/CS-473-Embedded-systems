// lt24_qsys.v

// Generated using ACDS version 13.1 182 at 2014.06.20.18:10:54

`timescale 1 ps / 1 ps
module lt24_qsys (
		input  wire        clk_clk,                                          //                                       clk.clk
		input  wire        reset_reset_n,                                    //                                     reset.reset_n
		output wire        lcd_reset_n_export,                               //                               lcd_reset_n.export
		input  wire        touch_panel_pen_irq_n_external_connection_export, // touch_panel_pen_irq_n_external_connection.export
		input  wire        touch_panel_busy_external_connection_export,      //      touch_panel_busy_external_connection.export
		input  wire        touch_panel_spi_external_MISO,                    //                  touch_panel_spi_external.MISO
		output wire        touch_panel_spi_external_MOSI,                    //                                          .MOSI
		output wire        touch_panel_spi_external_SCLK,                    //                                          .SCLK
		output wire        touch_panel_spi_external_SS_n,                    //                                          .SS_n
		input  wire        altpll_0_areset_conduit_export,                   //                   altpll_0_areset_conduit.export
		output wire        altpll_0_locked_conduit_export,                   //                   altpll_0_locked_conduit.export
		output wire        altpll_0_phasedone_conduit_export,                //                altpll_0_phasedone_conduit.export
		input  wire [3:0]  key_external_connection_export,                   //                   key_external_connection.export
		output wire        lt24_controller_0_conduit_end_cs,                 //             lt24_controller_0_conduit_end.cs
		output wire        lt24_controller_0_conduit_end_rs,                 //                                          .rs
		output wire        lt24_controller_0_conduit_end_rd,                 //                                          .rd
		output wire        lt24_controller_0_conduit_end_wr,                 //                                          .wr
		output wire [15:0] lt24_controller_0_conduit_end_data                //                                          .data
	);

	wire         altpll_sys_c1_clk;                                             // altpll_sys:c1 -> [LCD_RESET_N:clk, LT24_Controller_0:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, jtag_uart:clk, key:clk, mm_interconnect_0:altpll_sys_c1_clk, onchip_memory:clk, rst_controller_001:clk, sysid_qsys:clock, timer:clk, touch_panel_busy:clk, touch_panel_pen_irq_n:clk, touch_panel_spi:clk]
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;            // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;           // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire  [31:0] mm_interconnect_0_lcd_reset_n_s1_writedata;                    // mm_interconnect_0:LCD_RESET_N_s1_writedata -> LCD_RESET_N:writedata
	wire   [1:0] mm_interconnect_0_lcd_reset_n_s1_address;                      // mm_interconnect_0:LCD_RESET_N_s1_address -> LCD_RESET_N:address
	wire         mm_interconnect_0_lcd_reset_n_s1_chipselect;                   // mm_interconnect_0:LCD_RESET_N_s1_chipselect -> LCD_RESET_N:chipselect
	wire         mm_interconnect_0_lcd_reset_n_s1_write;                        // mm_interconnect_0:LCD_RESET_N_s1_write -> LCD_RESET_N:write_n
	wire  [31:0] mm_interconnect_0_lcd_reset_n_s1_readdata;                     // LCD_RESET_N:readdata -> mm_interconnect_0:LCD_RESET_N_s1_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                     // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [20:0] nios2_qsys_instruction_master_address;                         // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                            // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                        // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                   // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                          // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                            // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                         // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                              // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                           // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                              // mm_interconnect_0:key_s1_address -> key:address
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                             // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                  // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire  [16:0] mm_interconnect_0_onchip_memory_s1_address;                    // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                 // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire         mm_interconnect_0_onchip_memory_s1_clken;                      // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s1_write;                      // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                   // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                 // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire   [1:0] mm_interconnect_0_touch_panel_busy_s1_address;                 // mm_interconnect_0:touch_panel_busy_s1_address -> touch_panel_busy:address
	wire  [31:0] mm_interconnect_0_touch_panel_busy_s1_readdata;                // touch_panel_busy:readdata -> mm_interconnect_0:touch_panel_busy_s1_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest;    // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;      // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;        // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_write;          // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_read;           // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;       // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess;    // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;     // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire         nios2_qsys_data_master_waitrequest;                            // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                              // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [20:0] nios2_qsys_data_master_address;                                // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire         nios2_qsys_data_master_write;                                  // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire         nios2_qsys_data_master_read;                                   // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire  [31:0] nios2_qsys_data_master_readdata;                               // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                            // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                          // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                             // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire  [31:0] mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata;  // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_writedata -> LT24_Controller_0:s_writedata
	wire   [0:0] mm_interconnect_0_lt24_controller_0_avalon_slave_0_address;    // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_address -> LT24_Controller_0:s_address
	wire         mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect; // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_chipselect -> LT24_Controller_0:s_chipselect_n
	wire         mm_interconnect_0_lt24_controller_0_avalon_slave_0_write;      // mm_interconnect_0:LT24_Controller_0_avalon_slave_0_write -> LT24_Controller_0:s_write_n
	wire  [31:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata;          // mm_interconnect_0:touch_panel_pen_irq_n_s1_writedata -> touch_panel_pen_irq_n:writedata
	wire   [1:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_address;            // mm_interconnect_0:touch_panel_pen_irq_n_s1_address -> touch_panel_pen_irq_n:address
	wire         mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect;         // mm_interconnect_0:touch_panel_pen_irq_n_s1_chipselect -> touch_panel_pen_irq_n:chipselect
	wire         mm_interconnect_0_touch_panel_pen_irq_n_s1_write;              // mm_interconnect_0:touch_panel_pen_irq_n_s1_write -> touch_panel_pen_irq_n:write_n
	wire  [31:0] mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata;           // touch_panel_pen_irq_n:readdata -> mm_interconnect_0:touch_panel_pen_irq_n_s1_readdata
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;              // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire   [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;                // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire         mm_interconnect_0_altpll_sys_pll_slave_write;                  // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire         mm_interconnect_0_altpll_sys_pll_slave_read;                   // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;               // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_writedata;  // mm_interconnect_0:touch_panel_spi_spi_control_port_writedata -> touch_panel_spi:data_from_cpu
	wire   [2:0] mm_interconnect_0_touch_panel_spi_spi_control_port_address;    // mm_interconnect_0:touch_panel_spi_spi_control_port_address -> touch_panel_spi:mem_addr
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect; // mm_interconnect_0:touch_panel_spi_spi_control_port_chipselect -> touch_panel_spi:spi_select
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_write;      // mm_interconnect_0:touch_panel_spi_spi_control_port_write -> touch_panel_spi:write_n
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_read;       // mm_interconnect_0:touch_panel_spi_spi_control_port_read -> touch_panel_spi:read_n
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_readdata;   // touch_panel_spi:data_to_cpu -> mm_interconnect_0:touch_panel_spi_spi_control_port_readdata
	wire  [31:0] nios2_qsys_d_irq_irq;                                          // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire         irq_mapper_receiver0_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                 // jtag_uart:av_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                      // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                             // timer:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                      // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                             // touch_panel_spi:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                      // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                             // touch_panel_pen_irq_n:irq -> irq_synchronizer_003:receiver_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [nios2_qsys:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_jtag_debug_module_reset_reset;                      // nios2_qsys:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [LCD_RESET_N:reset_n, LT24_Controller_0:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, jtag_uart:rst_n, key:reset_n, mm_interconnect_0:onchip_memory_reset1_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator_001:in_reset, sysid_qsys:reset_n, timer:reset_n, touch_panel_busy:reset_n, touch_panel_pen_irq_n:reset_n, touch_panel_spi:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                        // rst_controller_001:reset_req -> [onchip_memory:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> [altpll_sys:reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset]

	lt24_qsys_nios2_qsys nios2_qsys (
		.clk                                   (clk_clk),                                                    //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	lt24_qsys_jtag_uart jtag_uart (
		.clk            (altpll_sys_c1_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_receiver_irq)                              //               irq.irq
	);

	lt24_qsys_onchip_memory onchip_memory (
		.clk        (altpll_sys_c1_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)         //       .reset_req
	);

	lt24_qsys_LCD_RESET_N lcd_reset_n (
		.clk        (altpll_sys_c1_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_lcd_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lcd_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lcd_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lcd_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lcd_reset_n_s1_readdata),   //                    .readdata
		.out_port   (lcd_reset_n_export)                           // external_connection.export
	);

	lt24_qsys_timer timer (
		.clk        (altpll_sys_c1_clk),                     //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)      //   irq.irq
	);

	lt24_qsys_touch_panel_spi touch_panel_spi (
		.clk           (altpll_sys_c1_clk),                                             //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                           //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_touch_panel_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_touch_panel_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_synchronizer_002_receiver_irq),                             //              irq.irq
		.MISO          (touch_panel_spi_external_MISO),                                 //         external.export
		.MOSI          (touch_panel_spi_external_MOSI),                                 //                 .export
		.SCLK          (touch_panel_spi_external_SCLK),                                 //                 .export
		.SS_n          (touch_panel_spi_external_SS_n)                                  //                 .export
	);

	lt24_qsys_touch_panel_pen_irq_n touch_panel_pen_irq_n (
		.clk        (altpll_sys_c1_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_touch_panel_pen_irq_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_panel_pen_irq_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata),   //                    .readdata
		.in_port    (touch_panel_pen_irq_n_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_003_receiver_irq)                      //                 irq.irq
	);

	lt24_qsys_touch_panel_busy touch_panel_busy (
		.clk      (altpll_sys_c1_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_touch_panel_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touch_panel_busy_s1_readdata), //                    .readdata
		.in_port  (touch_panel_busy_external_connection_export)     // external_connection.export
	);

	lt24_qsys_altpll_sys altpll_sys (
		.clk       (clk_clk),                                          //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0        (),                                                 //                    c0.clk
		.c1        (altpll_sys_c1_clk),                                //                    c1.clk
		.areset    (altpll_0_areset_conduit_export),                   //        areset_conduit.export
		.locked    (altpll_0_locked_conduit_export),                   //        locked_conduit.export
		.phasedone (altpll_0_phasedone_conduit_export)                 //     phasedone_conduit.export
	);

	lt24_qsys_key key (
		.clk      (altpll_sys_c1_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	LT24_Controller lt24_controller_0 (
		.clk            (altpll_sys_c1_clk),                                              //          clock.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                            //          reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect_n
		.s_write_n      (~mm_interconnect_0_lt24_controller_0_avalon_slave_0_write),      //               .write_n
		.s_writedata    (mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata),   //               .writedata
		.s_address      (mm_interconnect_0_lt24_controller_0_avalon_slave_0_address),     //               .address
		.lt24_cs        (lt24_controller_0_conduit_end_cs),                               //    conduit_end.export
		.lt24_rs        (lt24_controller_0_conduit_end_rs),                               //               .export
		.lt24_rd        (lt24_controller_0_conduit_end_rd),                               //               .export
		.lt24_wr        (lt24_controller_0_conduit_end_wr),                               //               .export
		.lt24_data      (lt24_controller_0_conduit_end_data)                              //               .export
	);

	lt24_qsys_sysid_qsys sysid_qsys (
		.clock    (altpll_sys_c1_clk),                                   //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	lt24_qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c1_clk                                            (altpll_sys_c1_clk),                                             //                                          altpll_sys_c1.clk
		.clk_50_clk_clk                                               (clk_clk),                                                       //                                             clk_50_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                            // altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                //               nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.onchip_memory_reset1_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                            //             onchip_memory_reset1_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                               (nios2_qsys_data_master_address),                                //                                 nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest                           (nios2_qsys_data_master_waitrequest),                            //                                                       .waitrequest
		.nios2_qsys_data_master_byteenable                            (nios2_qsys_data_master_byteenable),                             //                                                       .byteenable
		.nios2_qsys_data_master_read                                  (nios2_qsys_data_master_read),                                   //                                                       .read
		.nios2_qsys_data_master_readdata                              (nios2_qsys_data_master_readdata),                               //                                                       .readdata
		.nios2_qsys_data_master_readdatavalid                         (nios2_qsys_data_master_readdatavalid),                          //                                                       .readdatavalid
		.nios2_qsys_data_master_write                                 (nios2_qsys_data_master_write),                                  //                                                       .write
		.nios2_qsys_data_master_writedata                             (nios2_qsys_data_master_writedata),                              //                                                       .writedata
		.nios2_qsys_data_master_debugaccess                           (nios2_qsys_data_master_debugaccess),                            //                                                       .debugaccess
		.nios2_qsys_instruction_master_address                        (nios2_qsys_instruction_master_address),                         //                          nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest                    (nios2_qsys_instruction_master_waitrequest),                     //                                                       .waitrequest
		.nios2_qsys_instruction_master_read                           (nios2_qsys_instruction_master_read),                            //                                                       .read
		.nios2_qsys_instruction_master_readdata                       (nios2_qsys_instruction_master_readdata),                        //                                                       .readdata
		.nios2_qsys_instruction_master_readdatavalid                  (nios2_qsys_instruction_master_readdatavalid),                   //                                                       .readdatavalid
		.altpll_sys_pll_slave_address                                 (mm_interconnect_0_altpll_sys_pll_slave_address),                //                                   altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                   (mm_interconnect_0_altpll_sys_pll_slave_write),                  //                                                       .write
		.altpll_sys_pll_slave_read                                    (mm_interconnect_0_altpll_sys_pll_slave_read),                   //                                                       .read
		.altpll_sys_pll_slave_readdata                                (mm_interconnect_0_altpll_sys_pll_slave_readdata),               //                                                       .readdata
		.altpll_sys_pll_slave_writedata                               (mm_interconnect_0_altpll_sys_pll_slave_writedata),              //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                                       .chipselect
		.key_s1_address                                               (mm_interconnect_0_key_s1_address),                              //                                                 key_s1.address
		.key_s1_readdata                                              (mm_interconnect_0_key_s1_readdata),                             //                                                       .readdata
		.LCD_RESET_N_s1_address                                       (mm_interconnect_0_lcd_reset_n_s1_address),                      //                                         LCD_RESET_N_s1.address
		.LCD_RESET_N_s1_write                                         (mm_interconnect_0_lcd_reset_n_s1_write),                        //                                                       .write
		.LCD_RESET_N_s1_readdata                                      (mm_interconnect_0_lcd_reset_n_s1_readdata),                     //                                                       .readdata
		.LCD_RESET_N_s1_writedata                                     (mm_interconnect_0_lcd_reset_n_s1_writedata),                    //                                                       .writedata
		.LCD_RESET_N_s1_chipselect                                    (mm_interconnect_0_lcd_reset_n_s1_chipselect),                   //                                                       .chipselect
		.LT24_Controller_0_avalon_slave_0_address                     (mm_interconnect_0_lt24_controller_0_avalon_slave_0_address),    //                       LT24_Controller_0_avalon_slave_0.address
		.LT24_Controller_0_avalon_slave_0_write                       (mm_interconnect_0_lt24_controller_0_avalon_slave_0_write),      //                                                       .write
		.LT24_Controller_0_avalon_slave_0_writedata                   (mm_interconnect_0_lt24_controller_0_avalon_slave_0_writedata),  //                                                       .writedata
		.LT24_Controller_0_avalon_slave_0_chipselect                  (mm_interconnect_0_lt24_controller_0_avalon_slave_0_chipselect), //                                                       .chipselect
		.nios2_qsys_jtag_debug_module_address                         (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),        //                           nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write                           (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),          //                                                       .write
		.nios2_qsys_jtag_debug_module_read                            (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),           //                                                       .read
		.nios2_qsys_jtag_debug_module_readdata                        (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),       //                                                       .readdata
		.nios2_qsys_jtag_debug_module_writedata                       (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),      //                                                       .writedata
		.nios2_qsys_jtag_debug_module_byteenable                      (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),     //                                                       .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest                     (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest),    //                                                       .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess                     (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess),    //                                                       .debugaccess
		.onchip_memory_s1_address                                     (mm_interconnect_0_onchip_memory_s1_address),                    //                                       onchip_memory_s1.address
		.onchip_memory_s1_write                                       (mm_interconnect_0_onchip_memory_s1_write),                      //                                                       .write
		.onchip_memory_s1_readdata                                    (mm_interconnect_0_onchip_memory_s1_readdata),                   //                                                       .readdata
		.onchip_memory_s1_writedata                                   (mm_interconnect_0_onchip_memory_s1_writedata),                  //                                                       .writedata
		.onchip_memory_s1_byteenable                                  (mm_interconnect_0_onchip_memory_s1_byteenable),                 //                                                       .byteenable
		.onchip_memory_s1_chipselect                                  (mm_interconnect_0_onchip_memory_s1_chipselect),                 //                                                       .chipselect
		.onchip_memory_s1_clken                                       (mm_interconnect_0_onchip_memory_s1_clken),                      //                                                       .clken
		.sysid_qsys_control_slave_address                             (mm_interconnect_0_sysid_qsys_control_slave_address),            //                               sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                            (mm_interconnect_0_sysid_qsys_control_slave_readdata),           //                                                       .readdata
		.timer_s1_address                                             (mm_interconnect_0_timer_s1_address),                            //                                               timer_s1.address
		.timer_s1_write                                               (mm_interconnect_0_timer_s1_write),                              //                                                       .write
		.timer_s1_readdata                                            (mm_interconnect_0_timer_s1_readdata),                           //                                                       .readdata
		.timer_s1_writedata                                           (mm_interconnect_0_timer_s1_writedata),                          //                                                       .writedata
		.timer_s1_chipselect                                          (mm_interconnect_0_timer_s1_chipselect),                         //                                                       .chipselect
		.touch_panel_busy_s1_address                                  (mm_interconnect_0_touch_panel_busy_s1_address),                 //                                    touch_panel_busy_s1.address
		.touch_panel_busy_s1_readdata                                 (mm_interconnect_0_touch_panel_busy_s1_readdata),                //                                                       .readdata
		.touch_panel_pen_irq_n_s1_address                             (mm_interconnect_0_touch_panel_pen_irq_n_s1_address),            //                               touch_panel_pen_irq_n_s1.address
		.touch_panel_pen_irq_n_s1_write                               (mm_interconnect_0_touch_panel_pen_irq_n_s1_write),              //                                                       .write
		.touch_panel_pen_irq_n_s1_readdata                            (mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata),           //                                                       .readdata
		.touch_panel_pen_irq_n_s1_writedata                           (mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata),          //                                                       .writedata
		.touch_panel_pen_irq_n_s1_chipselect                          (mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect),         //                                                       .chipselect
		.touch_panel_spi_spi_control_port_address                     (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //                       touch_panel_spi_spi_control_port.address
		.touch_panel_spi_spi_control_port_write                       (mm_interconnect_0_touch_panel_spi_spi_control_port_write),      //                                                       .write
		.touch_panel_spi_spi_control_port_read                        (mm_interconnect_0_touch_panel_spi_spi_control_port_read),       //                                                       .read
		.touch_panel_spi_spi_control_port_readdata                    (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                                                       .readdata
		.touch_panel_spi_spi_control_port_writedata                   (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  //                                                       .writedata
		.touch_panel_spi_spi_control_port_chipselect                  (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect)  //                                                       .chipselect
	);

	lt24_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (altpll_sys_c1_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
