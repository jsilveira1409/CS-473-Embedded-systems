
module system2 (
	clk_clk,
	to_led_readdata);	

	input		clk_clk;
	output	[71:0]	to_led_readdata;
endmodule
