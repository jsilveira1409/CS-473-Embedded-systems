
module system (
	clk_clk,
	daisy_0_conduit_end_name,
	reset_reset_n);	

	input		clk_clk;
	output		daisy_0_conduit_end_name;
	input		reset_reset_n;
endmodule
