
module system2 (
	clk_clk,
	daisyport_0_conduit_end_writeresponsevalid_n);	

	input		clk_clk;
	output		daisyport_0_conduit_end_writeresponsevalid_n;
endmodule
