
module system (
	clk_clk,
	daisy_0_conduit_end_name);	

	input		clk_clk;
	output		daisy_0_conduit_end_name;
endmodule
