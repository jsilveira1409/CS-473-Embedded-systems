
module system (
	clk_clk,
	reset_reset_n,
	daisyport_0_conduit_end_name);	

	input		clk_clk;
	input		reset_reset_n;
	output		daisyport_0_conduit_end_name;
endmodule
